magic
tech gf180mcuC
magscale 1 5
timestamp 1670058501
<< obsm1 >>
rect 34449 4607 278591 228689
<< metal2 >>
rect 4900 297780 5012 298500
rect 13132 297780 13244 298500
rect 21364 297780 21476 298500
rect 29596 297780 29708 298500
rect 37828 297780 37940 298500
rect 46060 297780 46172 298500
rect 54292 297780 54404 298500
rect 62524 297780 62636 298500
rect 70756 297780 70868 298500
rect 78988 297780 79100 298500
rect 87220 297780 87332 298500
rect 95452 297780 95564 298500
rect 103684 297780 103796 298500
rect 111916 297780 112028 298500
rect 120148 297780 120260 298500
rect 128380 297780 128492 298500
rect 136612 297780 136724 298500
rect 144844 297780 144956 298500
rect 153076 297780 153188 298500
rect 161308 297780 161420 298500
rect 169540 297780 169652 298500
rect 177772 297780 177884 298500
rect 186004 297780 186116 298500
rect 194236 297780 194348 298500
rect 202468 297780 202580 298500
rect 210700 297780 210812 298500
rect 218932 297780 219044 298500
rect 227164 297780 227276 298500
rect 235396 297780 235508 298500
rect 243628 297780 243740 298500
rect 251860 297780 251972 298500
rect 260092 297780 260204 298500
rect 268324 297780 268436 298500
rect 276556 297780 276668 298500
rect 284788 297780 284900 298500
rect 293020 297780 293132 298500
rect 10892 -480 11004 240
rect 11452 -480 11564 240
rect 12012 -480 12124 240
rect 12572 -480 12684 240
rect 13132 -480 13244 240
rect 13692 -480 13804 240
rect 14252 -480 14364 240
rect 14812 -480 14924 240
rect 15372 -480 15484 240
rect 15932 -480 16044 240
rect 16492 -480 16604 240
rect 17052 -480 17164 240
rect 17612 -480 17724 240
rect 18172 -480 18284 240
rect 18732 -480 18844 240
rect 19292 -480 19404 240
rect 19852 -480 19964 240
rect 20412 -480 20524 240
rect 20972 -480 21084 240
rect 21532 -480 21644 240
rect 22092 -480 22204 240
rect 22652 -480 22764 240
rect 23212 -480 23324 240
rect 23772 -480 23884 240
rect 24332 -480 24444 240
rect 24892 -480 25004 240
rect 25452 -480 25564 240
rect 26012 -480 26124 240
rect 26572 -480 26684 240
rect 27132 -480 27244 240
rect 27692 -480 27804 240
rect 28252 -480 28364 240
rect 28812 -480 28924 240
rect 29372 -480 29484 240
rect 29932 -480 30044 240
rect 30492 -480 30604 240
rect 31052 -480 31164 240
rect 31612 -480 31724 240
rect 32172 -480 32284 240
rect 32732 -480 32844 240
rect 33292 -480 33404 240
rect 33852 -480 33964 240
rect 34412 -480 34524 240
rect 34972 -480 35084 240
rect 35532 -480 35644 240
rect 36092 -480 36204 240
rect 36652 -480 36764 240
rect 37212 -480 37324 240
rect 37772 -480 37884 240
rect 38332 -480 38444 240
rect 38892 -480 39004 240
rect 39452 -480 39564 240
rect 40012 -480 40124 240
rect 40572 -480 40684 240
rect 41132 -480 41244 240
rect 41692 -480 41804 240
rect 42252 -480 42364 240
rect 42812 -480 42924 240
rect 43372 -480 43484 240
rect 43932 -480 44044 240
rect 44492 -480 44604 240
rect 45052 -480 45164 240
rect 45612 -480 45724 240
rect 46172 -480 46284 240
rect 46732 -480 46844 240
rect 47292 -480 47404 240
rect 47852 -480 47964 240
rect 48412 -480 48524 240
rect 48972 -480 49084 240
rect 49532 -480 49644 240
rect 50092 -480 50204 240
rect 50652 -480 50764 240
rect 51212 -480 51324 240
rect 51772 -480 51884 240
rect 52332 -480 52444 240
rect 52892 -480 53004 240
rect 53452 -480 53564 240
rect 54012 -480 54124 240
rect 54572 -480 54684 240
rect 55132 -480 55244 240
rect 55692 -480 55804 240
rect 56252 -480 56364 240
rect 56812 -480 56924 240
rect 57372 -480 57484 240
rect 57932 -480 58044 240
rect 58492 -480 58604 240
rect 59052 -480 59164 240
rect 59612 -480 59724 240
rect 60172 -480 60284 240
rect 60732 -480 60844 240
rect 61292 -480 61404 240
rect 61852 -480 61964 240
rect 62412 -480 62524 240
rect 62972 -480 63084 240
rect 63532 -480 63644 240
rect 64092 -480 64204 240
rect 64652 -480 64764 240
rect 65212 -480 65324 240
rect 65772 -480 65884 240
rect 66332 -480 66444 240
rect 66892 -480 67004 240
rect 67452 -480 67564 240
rect 68012 -480 68124 240
rect 68572 -480 68684 240
rect 69132 -480 69244 240
rect 69692 -480 69804 240
rect 70252 -480 70364 240
rect 70812 -480 70924 240
rect 71372 -480 71484 240
rect 71932 -480 72044 240
rect 72492 -480 72604 240
rect 73052 -480 73164 240
rect 73612 -480 73724 240
rect 74172 -480 74284 240
rect 74732 -480 74844 240
rect 75292 -480 75404 240
rect 75852 -480 75964 240
rect 76412 -480 76524 240
rect 76972 -480 77084 240
rect 77532 -480 77644 240
rect 78092 -480 78204 240
rect 78652 -480 78764 240
rect 79212 -480 79324 240
rect 79772 -480 79884 240
rect 80332 -480 80444 240
rect 80892 -480 81004 240
rect 81452 -480 81564 240
rect 82012 -480 82124 240
rect 82572 -480 82684 240
rect 83132 -480 83244 240
rect 83692 -480 83804 240
rect 84252 -480 84364 240
rect 84812 -480 84924 240
rect 85372 -480 85484 240
rect 85932 -480 86044 240
rect 86492 -480 86604 240
rect 87052 -480 87164 240
rect 87612 -480 87724 240
rect 88172 -480 88284 240
rect 88732 -480 88844 240
rect 89292 -480 89404 240
rect 89852 -480 89964 240
rect 90412 -480 90524 240
rect 90972 -480 91084 240
rect 91532 -480 91644 240
rect 92092 -480 92204 240
rect 92652 -480 92764 240
rect 93212 -480 93324 240
rect 93772 -480 93884 240
rect 94332 -480 94444 240
rect 94892 -480 95004 240
rect 95452 -480 95564 240
rect 96012 -480 96124 240
rect 96572 -480 96684 240
rect 97132 -480 97244 240
rect 97692 -480 97804 240
rect 98252 -480 98364 240
rect 98812 -480 98924 240
rect 99372 -480 99484 240
rect 99932 -480 100044 240
rect 100492 -480 100604 240
rect 101052 -480 101164 240
rect 101612 -480 101724 240
rect 102172 -480 102284 240
rect 102732 -480 102844 240
rect 103292 -480 103404 240
rect 103852 -480 103964 240
rect 104412 -480 104524 240
rect 104972 -480 105084 240
rect 105532 -480 105644 240
rect 106092 -480 106204 240
rect 106652 -480 106764 240
rect 107212 -480 107324 240
rect 107772 -480 107884 240
rect 108332 -480 108444 240
rect 108892 -480 109004 240
rect 109452 -480 109564 240
rect 110012 -480 110124 240
rect 110572 -480 110684 240
rect 111132 -480 111244 240
rect 111692 -480 111804 240
rect 112252 -480 112364 240
rect 112812 -480 112924 240
rect 113372 -480 113484 240
rect 113932 -480 114044 240
rect 114492 -480 114604 240
rect 115052 -480 115164 240
rect 115612 -480 115724 240
rect 116172 -480 116284 240
rect 116732 -480 116844 240
rect 117292 -480 117404 240
rect 117852 -480 117964 240
rect 118412 -480 118524 240
rect 118972 -480 119084 240
rect 119532 -480 119644 240
rect 120092 -480 120204 240
rect 120652 -480 120764 240
rect 121212 -480 121324 240
rect 121772 -480 121884 240
rect 122332 -480 122444 240
rect 122892 -480 123004 240
rect 123452 -480 123564 240
rect 124012 -480 124124 240
rect 124572 -480 124684 240
rect 125132 -480 125244 240
rect 125692 -480 125804 240
rect 126252 -480 126364 240
rect 126812 -480 126924 240
rect 127372 -480 127484 240
rect 127932 -480 128044 240
rect 128492 -480 128604 240
rect 129052 -480 129164 240
rect 129612 -480 129724 240
rect 130172 -480 130284 240
rect 130732 -480 130844 240
rect 131292 -480 131404 240
rect 131852 -480 131964 240
rect 132412 -480 132524 240
rect 132972 -480 133084 240
rect 133532 -480 133644 240
rect 134092 -480 134204 240
rect 134652 -480 134764 240
rect 135212 -480 135324 240
rect 135772 -480 135884 240
rect 136332 -480 136444 240
rect 136892 -480 137004 240
rect 137452 -480 137564 240
rect 138012 -480 138124 240
rect 138572 -480 138684 240
rect 139132 -480 139244 240
rect 139692 -480 139804 240
rect 140252 -480 140364 240
rect 140812 -480 140924 240
rect 141372 -480 141484 240
rect 141932 -480 142044 240
rect 142492 -480 142604 240
rect 143052 -480 143164 240
rect 143612 -480 143724 240
rect 144172 -480 144284 240
rect 144732 -480 144844 240
rect 145292 -480 145404 240
rect 145852 -480 145964 240
rect 146412 -480 146524 240
rect 146972 -480 147084 240
rect 147532 -480 147644 240
rect 148092 -480 148204 240
rect 148652 -480 148764 240
rect 149212 -480 149324 240
rect 149772 -480 149884 240
rect 150332 -480 150444 240
rect 150892 -480 151004 240
rect 151452 -480 151564 240
rect 152012 -480 152124 240
rect 152572 -480 152684 240
rect 153132 -480 153244 240
rect 153692 -480 153804 240
rect 154252 -480 154364 240
rect 154812 -480 154924 240
rect 155372 -480 155484 240
rect 155932 -480 156044 240
rect 156492 -480 156604 240
rect 157052 -480 157164 240
rect 157612 -480 157724 240
rect 158172 -480 158284 240
rect 158732 -480 158844 240
rect 159292 -480 159404 240
rect 159852 -480 159964 240
rect 160412 -480 160524 240
rect 160972 -480 161084 240
rect 161532 -480 161644 240
rect 162092 -480 162204 240
rect 162652 -480 162764 240
rect 163212 -480 163324 240
rect 163772 -480 163884 240
rect 164332 -480 164444 240
rect 164892 -480 165004 240
rect 165452 -480 165564 240
rect 166012 -480 166124 240
rect 166572 -480 166684 240
rect 167132 -480 167244 240
rect 167692 -480 167804 240
rect 168252 -480 168364 240
rect 168812 -480 168924 240
rect 169372 -480 169484 240
rect 169932 -480 170044 240
rect 170492 -480 170604 240
rect 171052 -480 171164 240
rect 171612 -480 171724 240
rect 172172 -480 172284 240
rect 172732 -480 172844 240
rect 173292 -480 173404 240
rect 173852 -480 173964 240
rect 174412 -480 174524 240
rect 174972 -480 175084 240
rect 175532 -480 175644 240
rect 176092 -480 176204 240
rect 176652 -480 176764 240
rect 177212 -480 177324 240
rect 177772 -480 177884 240
rect 178332 -480 178444 240
rect 178892 -480 179004 240
rect 179452 -480 179564 240
rect 180012 -480 180124 240
rect 180572 -480 180684 240
rect 181132 -480 181244 240
rect 181692 -480 181804 240
rect 182252 -480 182364 240
rect 182812 -480 182924 240
rect 183372 -480 183484 240
rect 183932 -480 184044 240
rect 184492 -480 184604 240
rect 185052 -480 185164 240
rect 185612 -480 185724 240
rect 186172 -480 186284 240
rect 186732 -480 186844 240
rect 187292 -480 187404 240
rect 187852 -480 187964 240
rect 188412 -480 188524 240
rect 188972 -480 189084 240
rect 189532 -480 189644 240
rect 190092 -480 190204 240
rect 190652 -480 190764 240
rect 191212 -480 191324 240
rect 191772 -480 191884 240
rect 192332 -480 192444 240
rect 192892 -480 193004 240
rect 193452 -480 193564 240
rect 194012 -480 194124 240
rect 194572 -480 194684 240
rect 195132 -480 195244 240
rect 195692 -480 195804 240
rect 196252 -480 196364 240
rect 196812 -480 196924 240
rect 197372 -480 197484 240
rect 197932 -480 198044 240
rect 198492 -480 198604 240
rect 199052 -480 199164 240
rect 199612 -480 199724 240
rect 200172 -480 200284 240
rect 200732 -480 200844 240
rect 201292 -480 201404 240
rect 201852 -480 201964 240
rect 202412 -480 202524 240
rect 202972 -480 203084 240
rect 203532 -480 203644 240
rect 204092 -480 204204 240
rect 204652 -480 204764 240
rect 205212 -480 205324 240
rect 205772 -480 205884 240
rect 206332 -480 206444 240
rect 206892 -480 207004 240
rect 207452 -480 207564 240
rect 208012 -480 208124 240
rect 208572 -480 208684 240
rect 209132 -480 209244 240
rect 209692 -480 209804 240
rect 210252 -480 210364 240
rect 210812 -480 210924 240
rect 211372 -480 211484 240
rect 211932 -480 212044 240
rect 212492 -480 212604 240
rect 213052 -480 213164 240
rect 213612 -480 213724 240
rect 214172 -480 214284 240
rect 214732 -480 214844 240
rect 215292 -480 215404 240
rect 215852 -480 215964 240
rect 216412 -480 216524 240
rect 216972 -480 217084 240
rect 217532 -480 217644 240
rect 218092 -480 218204 240
rect 218652 -480 218764 240
rect 219212 -480 219324 240
rect 219772 -480 219884 240
rect 220332 -480 220444 240
rect 220892 -480 221004 240
rect 221452 -480 221564 240
rect 222012 -480 222124 240
rect 222572 -480 222684 240
rect 223132 -480 223244 240
rect 223692 -480 223804 240
rect 224252 -480 224364 240
rect 224812 -480 224924 240
rect 225372 -480 225484 240
rect 225932 -480 226044 240
rect 226492 -480 226604 240
rect 227052 -480 227164 240
rect 227612 -480 227724 240
rect 228172 -480 228284 240
rect 228732 -480 228844 240
rect 229292 -480 229404 240
rect 229852 -480 229964 240
rect 230412 -480 230524 240
rect 230972 -480 231084 240
rect 231532 -480 231644 240
rect 232092 -480 232204 240
rect 232652 -480 232764 240
rect 233212 -480 233324 240
rect 233772 -480 233884 240
rect 234332 -480 234444 240
rect 234892 -480 235004 240
rect 235452 -480 235564 240
rect 236012 -480 236124 240
rect 236572 -480 236684 240
rect 237132 -480 237244 240
rect 237692 -480 237804 240
rect 238252 -480 238364 240
rect 238812 -480 238924 240
rect 239372 -480 239484 240
rect 239932 -480 240044 240
rect 240492 -480 240604 240
rect 241052 -480 241164 240
rect 241612 -480 241724 240
rect 242172 -480 242284 240
rect 242732 -480 242844 240
rect 243292 -480 243404 240
rect 243852 -480 243964 240
rect 244412 -480 244524 240
rect 244972 -480 245084 240
rect 245532 -480 245644 240
rect 246092 -480 246204 240
rect 246652 -480 246764 240
rect 247212 -480 247324 240
rect 247772 -480 247884 240
rect 248332 -480 248444 240
rect 248892 -480 249004 240
rect 249452 -480 249564 240
rect 250012 -480 250124 240
rect 250572 -480 250684 240
rect 251132 -480 251244 240
rect 251692 -480 251804 240
rect 252252 -480 252364 240
rect 252812 -480 252924 240
rect 253372 -480 253484 240
rect 253932 -480 254044 240
rect 254492 -480 254604 240
rect 255052 -480 255164 240
rect 255612 -480 255724 240
rect 256172 -480 256284 240
rect 256732 -480 256844 240
rect 257292 -480 257404 240
rect 257852 -480 257964 240
rect 258412 -480 258524 240
rect 258972 -480 259084 240
rect 259532 -480 259644 240
rect 260092 -480 260204 240
rect 260652 -480 260764 240
rect 261212 -480 261324 240
rect 261772 -480 261884 240
rect 262332 -480 262444 240
rect 262892 -480 263004 240
rect 263452 -480 263564 240
rect 264012 -480 264124 240
rect 264572 -480 264684 240
rect 265132 -480 265244 240
rect 265692 -480 265804 240
rect 266252 -480 266364 240
rect 266812 -480 266924 240
rect 267372 -480 267484 240
rect 267932 -480 268044 240
rect 268492 -480 268604 240
rect 269052 -480 269164 240
rect 269612 -480 269724 240
rect 270172 -480 270284 240
rect 270732 -480 270844 240
rect 271292 -480 271404 240
rect 271852 -480 271964 240
rect 272412 -480 272524 240
rect 272972 -480 273084 240
rect 273532 -480 273644 240
rect 274092 -480 274204 240
rect 274652 -480 274764 240
rect 275212 -480 275324 240
rect 275772 -480 275884 240
rect 276332 -480 276444 240
rect 276892 -480 277004 240
rect 277452 -480 277564 240
rect 278012 -480 278124 240
rect 278572 -480 278684 240
rect 279132 -480 279244 240
rect 279692 -480 279804 240
rect 280252 -480 280364 240
rect 280812 -480 280924 240
rect 281372 -480 281484 240
rect 281932 -480 282044 240
rect 282492 -480 282604 240
rect 283052 -480 283164 240
rect 283612 -480 283724 240
rect 284172 -480 284284 240
rect 284732 -480 284844 240
rect 285292 -480 285404 240
rect 285852 -480 285964 240
rect 286412 -480 286524 240
rect 286972 -480 287084 240
<< obsm2 >>
rect 1246 297750 4870 297850
rect 5042 297750 13102 297850
rect 13274 297750 21334 297850
rect 21506 297750 29566 297850
rect 29738 297750 37798 297850
rect 37970 297750 46030 297850
rect 46202 297750 54262 297850
rect 54434 297750 62494 297850
rect 62666 297750 70726 297850
rect 70898 297750 78958 297850
rect 79130 297750 87190 297850
rect 87362 297750 95422 297850
rect 95594 297750 103654 297850
rect 103826 297750 111886 297850
rect 112058 297750 120118 297850
rect 120290 297750 128350 297850
rect 128522 297750 136582 297850
rect 136754 297750 144814 297850
rect 144986 297750 153046 297850
rect 153218 297750 161278 297850
rect 161450 297750 169510 297850
rect 169682 297750 177742 297850
rect 177914 297750 185974 297850
rect 186146 297750 194206 297850
rect 194378 297750 202438 297850
rect 202610 297750 210670 297850
rect 210842 297750 218902 297850
rect 219074 297750 227134 297850
rect 227306 297750 235366 297850
rect 235538 297750 243598 297850
rect 243770 297750 251830 297850
rect 252002 297750 260062 297850
rect 260234 297750 268294 297850
rect 268466 297750 276526 297850
rect 276698 297750 284758 297850
rect 284930 297750 292990 297850
rect 293162 297750 297010 297850
rect 1246 270 297010 297750
rect 1246 182 10862 270
rect 11034 182 11422 270
rect 11594 182 11982 270
rect 12154 182 12542 270
rect 12714 182 13102 270
rect 13274 182 13662 270
rect 13834 182 14222 270
rect 14394 182 14782 270
rect 14954 182 15342 270
rect 15514 182 15902 270
rect 16074 182 16462 270
rect 16634 182 17022 270
rect 17194 182 17582 270
rect 17754 182 18142 270
rect 18314 182 18702 270
rect 18874 182 19262 270
rect 19434 182 19822 270
rect 19994 182 20382 270
rect 20554 182 20942 270
rect 21114 182 21502 270
rect 21674 182 22062 270
rect 22234 182 22622 270
rect 22794 182 23182 270
rect 23354 182 23742 270
rect 23914 182 24302 270
rect 24474 182 24862 270
rect 25034 182 25422 270
rect 25594 182 25982 270
rect 26154 182 26542 270
rect 26714 182 27102 270
rect 27274 182 27662 270
rect 27834 182 28222 270
rect 28394 182 28782 270
rect 28954 182 29342 270
rect 29514 182 29902 270
rect 30074 182 30462 270
rect 30634 182 31022 270
rect 31194 182 31582 270
rect 31754 182 32142 270
rect 32314 182 32702 270
rect 32874 182 33262 270
rect 33434 182 33822 270
rect 33994 182 34382 270
rect 34554 182 34942 270
rect 35114 182 35502 270
rect 35674 182 36062 270
rect 36234 182 36622 270
rect 36794 182 37182 270
rect 37354 182 37742 270
rect 37914 182 38302 270
rect 38474 182 38862 270
rect 39034 182 39422 270
rect 39594 182 39982 270
rect 40154 182 40542 270
rect 40714 182 41102 270
rect 41274 182 41662 270
rect 41834 182 42222 270
rect 42394 182 42782 270
rect 42954 182 43342 270
rect 43514 182 43902 270
rect 44074 182 44462 270
rect 44634 182 45022 270
rect 45194 182 45582 270
rect 45754 182 46142 270
rect 46314 182 46702 270
rect 46874 182 47262 270
rect 47434 182 47822 270
rect 47994 182 48382 270
rect 48554 182 48942 270
rect 49114 182 49502 270
rect 49674 182 50062 270
rect 50234 182 50622 270
rect 50794 182 51182 270
rect 51354 182 51742 270
rect 51914 182 52302 270
rect 52474 182 52862 270
rect 53034 182 53422 270
rect 53594 182 53982 270
rect 54154 182 54542 270
rect 54714 182 55102 270
rect 55274 182 55662 270
rect 55834 182 56222 270
rect 56394 182 56782 270
rect 56954 182 57342 270
rect 57514 182 57902 270
rect 58074 182 58462 270
rect 58634 182 59022 270
rect 59194 182 59582 270
rect 59754 182 60142 270
rect 60314 182 60702 270
rect 60874 182 61262 270
rect 61434 182 61822 270
rect 61994 182 62382 270
rect 62554 182 62942 270
rect 63114 182 63502 270
rect 63674 182 64062 270
rect 64234 182 64622 270
rect 64794 182 65182 270
rect 65354 182 65742 270
rect 65914 182 66302 270
rect 66474 182 66862 270
rect 67034 182 67422 270
rect 67594 182 67982 270
rect 68154 182 68542 270
rect 68714 182 69102 270
rect 69274 182 69662 270
rect 69834 182 70222 270
rect 70394 182 70782 270
rect 70954 182 71342 270
rect 71514 182 71902 270
rect 72074 182 72462 270
rect 72634 182 73022 270
rect 73194 182 73582 270
rect 73754 182 74142 270
rect 74314 182 74702 270
rect 74874 182 75262 270
rect 75434 182 75822 270
rect 75994 182 76382 270
rect 76554 182 76942 270
rect 77114 182 77502 270
rect 77674 182 78062 270
rect 78234 182 78622 270
rect 78794 182 79182 270
rect 79354 182 79742 270
rect 79914 182 80302 270
rect 80474 182 80862 270
rect 81034 182 81422 270
rect 81594 182 81982 270
rect 82154 182 82542 270
rect 82714 182 83102 270
rect 83274 182 83662 270
rect 83834 182 84222 270
rect 84394 182 84782 270
rect 84954 182 85342 270
rect 85514 182 85902 270
rect 86074 182 86462 270
rect 86634 182 87022 270
rect 87194 182 87582 270
rect 87754 182 88142 270
rect 88314 182 88702 270
rect 88874 182 89262 270
rect 89434 182 89822 270
rect 89994 182 90382 270
rect 90554 182 90942 270
rect 91114 182 91502 270
rect 91674 182 92062 270
rect 92234 182 92622 270
rect 92794 182 93182 270
rect 93354 182 93742 270
rect 93914 182 94302 270
rect 94474 182 94862 270
rect 95034 182 95422 270
rect 95594 182 95982 270
rect 96154 182 96542 270
rect 96714 182 97102 270
rect 97274 182 97662 270
rect 97834 182 98222 270
rect 98394 182 98782 270
rect 98954 182 99342 270
rect 99514 182 99902 270
rect 100074 182 100462 270
rect 100634 182 101022 270
rect 101194 182 101582 270
rect 101754 182 102142 270
rect 102314 182 102702 270
rect 102874 182 103262 270
rect 103434 182 103822 270
rect 103994 182 104382 270
rect 104554 182 104942 270
rect 105114 182 105502 270
rect 105674 182 106062 270
rect 106234 182 106622 270
rect 106794 182 107182 270
rect 107354 182 107742 270
rect 107914 182 108302 270
rect 108474 182 108862 270
rect 109034 182 109422 270
rect 109594 182 109982 270
rect 110154 182 110542 270
rect 110714 182 111102 270
rect 111274 182 111662 270
rect 111834 182 112222 270
rect 112394 182 112782 270
rect 112954 182 113342 270
rect 113514 182 113902 270
rect 114074 182 114462 270
rect 114634 182 115022 270
rect 115194 182 115582 270
rect 115754 182 116142 270
rect 116314 182 116702 270
rect 116874 182 117262 270
rect 117434 182 117822 270
rect 117994 182 118382 270
rect 118554 182 118942 270
rect 119114 182 119502 270
rect 119674 182 120062 270
rect 120234 182 120622 270
rect 120794 182 121182 270
rect 121354 182 121742 270
rect 121914 182 122302 270
rect 122474 182 122862 270
rect 123034 182 123422 270
rect 123594 182 123982 270
rect 124154 182 124542 270
rect 124714 182 125102 270
rect 125274 182 125662 270
rect 125834 182 126222 270
rect 126394 182 126782 270
rect 126954 182 127342 270
rect 127514 182 127902 270
rect 128074 182 128462 270
rect 128634 182 129022 270
rect 129194 182 129582 270
rect 129754 182 130142 270
rect 130314 182 130702 270
rect 130874 182 131262 270
rect 131434 182 131822 270
rect 131994 182 132382 270
rect 132554 182 132942 270
rect 133114 182 133502 270
rect 133674 182 134062 270
rect 134234 182 134622 270
rect 134794 182 135182 270
rect 135354 182 135742 270
rect 135914 182 136302 270
rect 136474 182 136862 270
rect 137034 182 137422 270
rect 137594 182 137982 270
rect 138154 182 138542 270
rect 138714 182 139102 270
rect 139274 182 139662 270
rect 139834 182 140222 270
rect 140394 182 140782 270
rect 140954 182 141342 270
rect 141514 182 141902 270
rect 142074 182 142462 270
rect 142634 182 143022 270
rect 143194 182 143582 270
rect 143754 182 144142 270
rect 144314 182 144702 270
rect 144874 182 145262 270
rect 145434 182 145822 270
rect 145994 182 146382 270
rect 146554 182 146942 270
rect 147114 182 147502 270
rect 147674 182 148062 270
rect 148234 182 148622 270
rect 148794 182 149182 270
rect 149354 182 149742 270
rect 149914 182 150302 270
rect 150474 182 150862 270
rect 151034 182 151422 270
rect 151594 182 151982 270
rect 152154 182 152542 270
rect 152714 182 153102 270
rect 153274 182 153662 270
rect 153834 182 154222 270
rect 154394 182 154782 270
rect 154954 182 155342 270
rect 155514 182 155902 270
rect 156074 182 156462 270
rect 156634 182 157022 270
rect 157194 182 157582 270
rect 157754 182 158142 270
rect 158314 182 158702 270
rect 158874 182 159262 270
rect 159434 182 159822 270
rect 159994 182 160382 270
rect 160554 182 160942 270
rect 161114 182 161502 270
rect 161674 182 162062 270
rect 162234 182 162622 270
rect 162794 182 163182 270
rect 163354 182 163742 270
rect 163914 182 164302 270
rect 164474 182 164862 270
rect 165034 182 165422 270
rect 165594 182 165982 270
rect 166154 182 166542 270
rect 166714 182 167102 270
rect 167274 182 167662 270
rect 167834 182 168222 270
rect 168394 182 168782 270
rect 168954 182 169342 270
rect 169514 182 169902 270
rect 170074 182 170462 270
rect 170634 182 171022 270
rect 171194 182 171582 270
rect 171754 182 172142 270
rect 172314 182 172702 270
rect 172874 182 173262 270
rect 173434 182 173822 270
rect 173994 182 174382 270
rect 174554 182 174942 270
rect 175114 182 175502 270
rect 175674 182 176062 270
rect 176234 182 176622 270
rect 176794 182 177182 270
rect 177354 182 177742 270
rect 177914 182 178302 270
rect 178474 182 178862 270
rect 179034 182 179422 270
rect 179594 182 179982 270
rect 180154 182 180542 270
rect 180714 182 181102 270
rect 181274 182 181662 270
rect 181834 182 182222 270
rect 182394 182 182782 270
rect 182954 182 183342 270
rect 183514 182 183902 270
rect 184074 182 184462 270
rect 184634 182 185022 270
rect 185194 182 185582 270
rect 185754 182 186142 270
rect 186314 182 186702 270
rect 186874 182 187262 270
rect 187434 182 187822 270
rect 187994 182 188382 270
rect 188554 182 188942 270
rect 189114 182 189502 270
rect 189674 182 190062 270
rect 190234 182 190622 270
rect 190794 182 191182 270
rect 191354 182 191742 270
rect 191914 182 192302 270
rect 192474 182 192862 270
rect 193034 182 193422 270
rect 193594 182 193982 270
rect 194154 182 194542 270
rect 194714 182 195102 270
rect 195274 182 195662 270
rect 195834 182 196222 270
rect 196394 182 196782 270
rect 196954 182 197342 270
rect 197514 182 197902 270
rect 198074 182 198462 270
rect 198634 182 199022 270
rect 199194 182 199582 270
rect 199754 182 200142 270
rect 200314 182 200702 270
rect 200874 182 201262 270
rect 201434 182 201822 270
rect 201994 182 202382 270
rect 202554 182 202942 270
rect 203114 182 203502 270
rect 203674 182 204062 270
rect 204234 182 204622 270
rect 204794 182 205182 270
rect 205354 182 205742 270
rect 205914 182 206302 270
rect 206474 182 206862 270
rect 207034 182 207422 270
rect 207594 182 207982 270
rect 208154 182 208542 270
rect 208714 182 209102 270
rect 209274 182 209662 270
rect 209834 182 210222 270
rect 210394 182 210782 270
rect 210954 182 211342 270
rect 211514 182 211902 270
rect 212074 182 212462 270
rect 212634 182 213022 270
rect 213194 182 213582 270
rect 213754 182 214142 270
rect 214314 182 214702 270
rect 214874 182 215262 270
rect 215434 182 215822 270
rect 215994 182 216382 270
rect 216554 182 216942 270
rect 217114 182 217502 270
rect 217674 182 218062 270
rect 218234 182 218622 270
rect 218794 182 219182 270
rect 219354 182 219742 270
rect 219914 182 220302 270
rect 220474 182 220862 270
rect 221034 182 221422 270
rect 221594 182 221982 270
rect 222154 182 222542 270
rect 222714 182 223102 270
rect 223274 182 223662 270
rect 223834 182 224222 270
rect 224394 182 224782 270
rect 224954 182 225342 270
rect 225514 182 225902 270
rect 226074 182 226462 270
rect 226634 182 227022 270
rect 227194 182 227582 270
rect 227754 182 228142 270
rect 228314 182 228702 270
rect 228874 182 229262 270
rect 229434 182 229822 270
rect 229994 182 230382 270
rect 230554 182 230942 270
rect 231114 182 231502 270
rect 231674 182 232062 270
rect 232234 182 232622 270
rect 232794 182 233182 270
rect 233354 182 233742 270
rect 233914 182 234302 270
rect 234474 182 234862 270
rect 235034 182 235422 270
rect 235594 182 235982 270
rect 236154 182 236542 270
rect 236714 182 237102 270
rect 237274 182 237662 270
rect 237834 182 238222 270
rect 238394 182 238782 270
rect 238954 182 239342 270
rect 239514 182 239902 270
rect 240074 182 240462 270
rect 240634 182 241022 270
rect 241194 182 241582 270
rect 241754 182 242142 270
rect 242314 182 242702 270
rect 242874 182 243262 270
rect 243434 182 243822 270
rect 243994 182 244382 270
rect 244554 182 244942 270
rect 245114 182 245502 270
rect 245674 182 246062 270
rect 246234 182 246622 270
rect 246794 182 247182 270
rect 247354 182 247742 270
rect 247914 182 248302 270
rect 248474 182 248862 270
rect 249034 182 249422 270
rect 249594 182 249982 270
rect 250154 182 250542 270
rect 250714 182 251102 270
rect 251274 182 251662 270
rect 251834 182 252222 270
rect 252394 182 252782 270
rect 252954 182 253342 270
rect 253514 182 253902 270
rect 254074 182 254462 270
rect 254634 182 255022 270
rect 255194 182 255582 270
rect 255754 182 256142 270
rect 256314 182 256702 270
rect 256874 182 257262 270
rect 257434 182 257822 270
rect 257994 182 258382 270
rect 258554 182 258942 270
rect 259114 182 259502 270
rect 259674 182 260062 270
rect 260234 182 260622 270
rect 260794 182 261182 270
rect 261354 182 261742 270
rect 261914 182 262302 270
rect 262474 182 262862 270
rect 263034 182 263422 270
rect 263594 182 263982 270
rect 264154 182 264542 270
rect 264714 182 265102 270
rect 265274 182 265662 270
rect 265834 182 266222 270
rect 266394 182 266782 270
rect 266954 182 267342 270
rect 267514 182 267902 270
rect 268074 182 268462 270
rect 268634 182 269022 270
rect 269194 182 269582 270
rect 269754 182 270142 270
rect 270314 182 270702 270
rect 270874 182 271262 270
rect 271434 182 271822 270
rect 271994 182 272382 270
rect 272554 182 272942 270
rect 273114 182 273502 270
rect 273674 182 274062 270
rect 274234 182 274622 270
rect 274794 182 275182 270
rect 275354 182 275742 270
rect 275914 182 276302 270
rect 276474 182 276862 270
rect 277034 182 277422 270
rect 277594 182 277982 270
rect 278154 182 278542 270
rect 278714 182 279102 270
rect 279274 182 279662 270
rect 279834 182 280222 270
rect 280394 182 280782 270
rect 280954 182 281342 270
rect 281514 182 281902 270
rect 282074 182 282462 270
rect 282634 182 283022 270
rect 283194 182 283582 270
rect 283754 182 284142 270
rect 284314 182 284702 270
rect 284874 182 285262 270
rect 285434 182 285822 270
rect 285994 182 286382 270
rect 286554 182 286942 270
rect 287114 182 297010 270
<< metal3 >>
rect 297780 294532 298500 294644
rect -480 294364 240 294476
rect -480 288876 240 288988
rect 297780 288932 298500 289044
rect -480 283388 240 283500
rect 297780 283332 298500 283444
rect -480 277900 240 278012
rect 297780 277732 298500 277844
rect -480 272412 240 272524
rect 297780 272132 298500 272244
rect -480 266924 240 267036
rect 297780 266532 298500 266644
rect -480 261436 240 261548
rect 297780 260932 298500 261044
rect -480 255948 240 256060
rect 297780 255332 298500 255444
rect -480 250460 240 250572
rect 297780 249732 298500 249844
rect -480 244972 240 245084
rect 297780 244132 298500 244244
rect -480 239484 240 239596
rect 297780 238532 298500 238644
rect -480 233996 240 234108
rect 297780 232932 298500 233044
rect -480 228508 240 228620
rect 297780 227332 298500 227444
rect -480 223020 240 223132
rect 297780 221732 298500 221844
rect -480 217532 240 217644
rect 297780 216132 298500 216244
rect -480 212044 240 212156
rect 297780 210532 298500 210644
rect -480 206556 240 206668
rect 297780 204932 298500 205044
rect -480 201068 240 201180
rect 297780 199332 298500 199444
rect -480 195580 240 195692
rect 297780 193732 298500 193844
rect -480 190092 240 190204
rect 297780 188132 298500 188244
rect -480 184604 240 184716
rect 297780 182532 298500 182644
rect -480 179116 240 179228
rect 297780 176932 298500 177044
rect -480 173628 240 173740
rect 297780 171332 298500 171444
rect -480 168140 240 168252
rect 297780 165732 298500 165844
rect -480 162652 240 162764
rect 297780 160132 298500 160244
rect -480 157164 240 157276
rect 297780 154532 298500 154644
rect -480 151676 240 151788
rect 297780 148932 298500 149044
rect -480 146188 240 146300
rect 297780 143332 298500 143444
rect -480 140700 240 140812
rect 297780 137732 298500 137844
rect -480 135212 240 135324
rect 297780 132132 298500 132244
rect -480 129724 240 129836
rect 297780 126532 298500 126644
rect -480 124236 240 124348
rect 297780 120932 298500 121044
rect -480 118748 240 118860
rect 297780 115332 298500 115444
rect -480 113260 240 113372
rect 297780 109732 298500 109844
rect -480 107772 240 107884
rect 297780 104132 298500 104244
rect -480 102284 240 102396
rect 297780 98532 298500 98644
rect -480 96796 240 96908
rect 297780 92932 298500 93044
rect -480 91308 240 91420
rect 297780 87332 298500 87444
rect -480 85820 240 85932
rect 297780 81732 298500 81844
rect -480 80332 240 80444
rect 297780 76132 298500 76244
rect -480 74844 240 74956
rect 297780 70532 298500 70644
rect -480 69356 240 69468
rect 297780 64932 298500 65044
rect -480 63868 240 63980
rect 297780 59332 298500 59444
rect -480 58380 240 58492
rect 297780 53732 298500 53844
rect -480 52892 240 53004
rect 297780 48132 298500 48244
rect -480 47404 240 47516
rect 297780 42532 298500 42644
rect -480 41916 240 42028
rect 297780 36932 298500 37044
rect -480 36428 240 36540
rect 297780 31332 298500 31444
rect -480 30940 240 31052
rect 297780 25732 298500 25844
rect -480 25452 240 25564
rect 297780 20132 298500 20244
rect -480 19964 240 20076
rect -480 14476 240 14588
rect 297780 14532 298500 14644
rect -480 8988 240 9100
rect 297780 8932 298500 9044
rect -480 3500 240 3612
rect 297780 3332 298500 3444
<< obsm3 >>
rect 182 294674 297850 295666
rect 182 294506 297750 294674
rect 270 294502 297750 294506
rect 270 294334 297850 294502
rect 182 289074 297850 294334
rect 182 289018 297750 289074
rect 270 288902 297750 289018
rect 270 288846 297850 288902
rect 182 283530 297850 288846
rect 270 283474 297850 283530
rect 270 283358 297750 283474
rect 182 283302 297750 283358
rect 182 278042 297850 283302
rect 270 277874 297850 278042
rect 270 277870 297750 277874
rect 182 277702 297750 277870
rect 182 272554 297850 277702
rect 270 272382 297850 272554
rect 182 272274 297850 272382
rect 182 272102 297750 272274
rect 182 267066 297850 272102
rect 270 266894 297850 267066
rect 182 266674 297850 266894
rect 182 266502 297750 266674
rect 182 261578 297850 266502
rect 270 261406 297850 261578
rect 182 261074 297850 261406
rect 182 260902 297750 261074
rect 182 256090 297850 260902
rect 270 255918 297850 256090
rect 182 255474 297850 255918
rect 182 255302 297750 255474
rect 182 250602 297850 255302
rect 270 250430 297850 250602
rect 182 249874 297850 250430
rect 182 249702 297750 249874
rect 182 245114 297850 249702
rect 270 244942 297850 245114
rect 182 244274 297850 244942
rect 182 244102 297750 244274
rect 182 239626 297850 244102
rect 270 239454 297850 239626
rect 182 238674 297850 239454
rect 182 238502 297750 238674
rect 182 234138 297850 238502
rect 270 233966 297850 234138
rect 182 233074 297850 233966
rect 182 232902 297750 233074
rect 182 228650 297850 232902
rect 270 228478 297850 228650
rect 182 227474 297850 228478
rect 182 227302 297750 227474
rect 182 223162 297850 227302
rect 270 222990 297850 223162
rect 182 221874 297850 222990
rect 182 221702 297750 221874
rect 182 217674 297850 221702
rect 270 217502 297850 217674
rect 182 216274 297850 217502
rect 182 216102 297750 216274
rect 182 212186 297850 216102
rect 270 212014 297850 212186
rect 182 210674 297850 212014
rect 182 210502 297750 210674
rect 182 206698 297850 210502
rect 270 206526 297850 206698
rect 182 205074 297850 206526
rect 182 204902 297750 205074
rect 182 201210 297850 204902
rect 270 201038 297850 201210
rect 182 199474 297850 201038
rect 182 199302 297750 199474
rect 182 195722 297850 199302
rect 270 195550 297850 195722
rect 182 193874 297850 195550
rect 182 193702 297750 193874
rect 182 190234 297850 193702
rect 270 190062 297850 190234
rect 182 188274 297850 190062
rect 182 188102 297750 188274
rect 182 184746 297850 188102
rect 270 184574 297850 184746
rect 182 182674 297850 184574
rect 182 182502 297750 182674
rect 182 179258 297850 182502
rect 270 179086 297850 179258
rect 182 177074 297850 179086
rect 182 176902 297750 177074
rect 182 173770 297850 176902
rect 270 173598 297850 173770
rect 182 171474 297850 173598
rect 182 171302 297750 171474
rect 182 168282 297850 171302
rect 270 168110 297850 168282
rect 182 165874 297850 168110
rect 182 165702 297750 165874
rect 182 162794 297850 165702
rect 270 162622 297850 162794
rect 182 160274 297850 162622
rect 182 160102 297750 160274
rect 182 157306 297850 160102
rect 270 157134 297850 157306
rect 182 154674 297850 157134
rect 182 154502 297750 154674
rect 182 151818 297850 154502
rect 270 151646 297850 151818
rect 182 149074 297850 151646
rect 182 148902 297750 149074
rect 182 146330 297850 148902
rect 270 146158 297850 146330
rect 182 143474 297850 146158
rect 182 143302 297750 143474
rect 182 140842 297850 143302
rect 270 140670 297850 140842
rect 182 137874 297850 140670
rect 182 137702 297750 137874
rect 182 135354 297850 137702
rect 270 135182 297850 135354
rect 182 132274 297850 135182
rect 182 132102 297750 132274
rect 182 129866 297850 132102
rect 270 129694 297850 129866
rect 182 126674 297850 129694
rect 182 126502 297750 126674
rect 182 124378 297850 126502
rect 270 124206 297850 124378
rect 182 121074 297850 124206
rect 182 120902 297750 121074
rect 182 118890 297850 120902
rect 270 118718 297850 118890
rect 182 115474 297850 118718
rect 182 115302 297750 115474
rect 182 113402 297850 115302
rect 270 113230 297850 113402
rect 182 109874 297850 113230
rect 182 109702 297750 109874
rect 182 107914 297850 109702
rect 270 107742 297850 107914
rect 182 104274 297850 107742
rect 182 104102 297750 104274
rect 182 102426 297850 104102
rect 270 102254 297850 102426
rect 182 98674 297850 102254
rect 182 98502 297750 98674
rect 182 96938 297850 98502
rect 270 96766 297850 96938
rect 182 93074 297850 96766
rect 182 92902 297750 93074
rect 182 91450 297850 92902
rect 270 91278 297850 91450
rect 182 87474 297850 91278
rect 182 87302 297750 87474
rect 182 85962 297850 87302
rect 270 85790 297850 85962
rect 182 81874 297850 85790
rect 182 81702 297750 81874
rect 182 80474 297850 81702
rect 270 80302 297850 80474
rect 182 76274 297850 80302
rect 182 76102 297750 76274
rect 182 74986 297850 76102
rect 270 74814 297850 74986
rect 182 70674 297850 74814
rect 182 70502 297750 70674
rect 182 69498 297850 70502
rect 270 69326 297850 69498
rect 182 65074 297850 69326
rect 182 64902 297750 65074
rect 182 64010 297850 64902
rect 270 63838 297850 64010
rect 182 59474 297850 63838
rect 182 59302 297750 59474
rect 182 58522 297850 59302
rect 270 58350 297850 58522
rect 182 53874 297850 58350
rect 182 53702 297750 53874
rect 182 53034 297850 53702
rect 270 52862 297850 53034
rect 182 48274 297850 52862
rect 182 48102 297750 48274
rect 182 47546 297850 48102
rect 270 47374 297850 47546
rect 182 42674 297850 47374
rect 182 42502 297750 42674
rect 182 42058 297850 42502
rect 270 41886 297850 42058
rect 182 37074 297850 41886
rect 182 36902 297750 37074
rect 182 36570 297850 36902
rect 270 36398 297850 36570
rect 182 31474 297850 36398
rect 182 31302 297750 31474
rect 182 31082 297850 31302
rect 270 30910 297850 31082
rect 182 25874 297850 30910
rect 182 25702 297750 25874
rect 182 25594 297850 25702
rect 270 25422 297850 25594
rect 182 20274 297850 25422
rect 182 20106 297750 20274
rect 270 20102 297750 20106
rect 270 19934 297850 20102
rect 182 14674 297850 19934
rect 182 14618 297750 14674
rect 270 14502 297750 14618
rect 270 14446 297850 14502
rect 182 9130 297850 14446
rect 270 9074 297850 9130
rect 270 8958 297750 9074
rect 182 8902 297750 8958
rect 182 3642 297850 8902
rect 270 3474 297850 3642
rect 270 3470 297750 3474
rect 182 3302 297750 3470
rect 182 1806 297850 3302
<< metal4 >>
rect -958 -822 -648 299134
rect -478 -342 -168 298654
rect 1577 -822 1887 299134
rect 3437 -822 3747 299134
rect 10577 -822 10887 299134
rect 12437 -822 12747 299134
rect 19577 -822 19887 299134
rect 21437 -822 21747 299134
rect 28577 -822 28887 299134
rect 30437 -822 30747 299134
rect 37577 -822 37887 299134
rect 39437 -822 39747 299134
rect 46577 -822 46887 299134
rect 48437 -822 48747 299134
rect 55577 -822 55887 299134
rect 57437 -822 57747 299134
rect 64577 -822 64887 299134
rect 66437 -822 66747 299134
rect 73577 -822 73887 299134
rect 75437 -822 75747 299134
rect 82577 -822 82887 299134
rect 84437 -822 84747 299134
rect 91577 -822 91887 299134
rect 93437 -822 93747 299134
rect 100577 -822 100887 299134
rect 102437 -822 102747 299134
rect 109577 -822 109887 299134
rect 111437 -822 111747 299134
rect 118577 -822 118887 299134
rect 120437 -822 120747 299134
rect 127577 228466 127887 299134
rect 127577 -822 127887 169510
rect 129437 -822 129747 299134
rect 136577 -822 136887 299134
rect 138437 -822 138747 299134
rect 145577 -822 145887 299134
rect 147437 -822 147747 299134
rect 154577 -822 154887 299134
rect 156437 -822 156747 299134
rect 163577 -822 163887 299134
rect 165437 -822 165747 299134
rect 172577 228091 172887 299134
rect 174437 228091 174747 299134
rect 172577 -822 172887 224765
rect 174437 -822 174747 224765
rect 181577 -822 181887 299134
rect 183437 -822 183747 299134
rect 190577 -822 190887 299134
rect 192437 -822 192747 299134
rect 199577 -822 199887 299134
rect 201437 -822 201747 299134
rect 208577 -822 208887 299134
rect 210437 -822 210747 299134
rect 217577 -822 217887 299134
rect 219437 -822 219747 299134
rect 226577 -822 226887 299134
rect 228437 -822 228747 299134
rect 235577 -822 235887 299134
rect 237437 -822 237747 299134
rect 244577 -822 244887 299134
rect 246437 -822 246747 299134
rect 253577 -822 253887 299134
rect 255437 -822 255747 299134
rect 262577 -822 262887 299134
rect 264437 -822 264747 299134
rect 271577 -822 271887 299134
rect 273437 -822 273747 299134
rect 280577 -822 280887 299134
rect 282437 -822 282747 299134
rect 289577 -822 289887 299134
rect 291437 -822 291747 299134
rect 298200 -342 298510 298654
rect 298680 -822 298990 299134
<< obsm4 >>
rect 36974 1969 37547 229815
rect 37917 1969 39407 229815
rect 39777 1969 46547 229815
rect 46917 1969 48407 229815
rect 48777 1969 55547 229815
rect 55917 1969 57407 229815
rect 57777 1969 64547 229815
rect 64917 1969 66407 229815
rect 66777 1969 73547 229815
rect 73917 1969 75407 229815
rect 75777 1969 82547 229815
rect 82917 1969 84407 229815
rect 84777 1969 91547 229815
rect 91917 1969 93407 229815
rect 93777 1969 100547 229815
rect 100917 1969 102407 229815
rect 102777 1969 109547 229815
rect 109917 1969 111407 229815
rect 111777 1969 118547 229815
rect 118917 1969 120407 229815
rect 120777 228436 127547 229815
rect 127917 228436 129407 229815
rect 120777 169540 129407 228436
rect 120777 1969 127547 169540
rect 127917 1969 129407 169540
rect 129777 1969 136547 229815
rect 136917 1969 138407 229815
rect 138777 1969 145547 229815
rect 145917 1969 147407 229815
rect 147777 1969 154547 229815
rect 154917 1969 156407 229815
rect 156777 1969 163547 229815
rect 163917 1969 165407 229815
rect 165777 228061 172547 229815
rect 172917 228061 174407 229815
rect 174777 228061 181547 229815
rect 165777 224795 181547 228061
rect 165777 1969 172547 224795
rect 172917 1969 174407 224795
rect 174777 1969 181547 224795
rect 181917 1969 183407 229815
rect 183777 1969 190547 229815
rect 190917 1969 192407 229815
rect 192777 1969 199547 229815
rect 199917 1969 201407 229815
rect 201777 1969 208547 229815
rect 208917 1969 210407 229815
rect 210777 1969 217547 229815
rect 217917 1969 219407 229815
rect 219777 1969 226547 229815
rect 226917 1969 228407 229815
rect 228777 1969 235547 229815
rect 235917 1969 237407 229815
rect 237777 1969 244547 229815
rect 244917 1969 246407 229815
rect 246777 1969 251314 229815
<< metal5 >>
rect -958 298824 298990 299134
rect -478 298344 298510 298654
rect -958 292913 298990 293223
rect -958 289913 298990 290223
rect -958 283913 298990 284223
rect -958 280913 298990 281223
rect -958 274913 298990 275223
rect -958 271913 298990 272223
rect -958 265913 298990 266223
rect -958 262913 298990 263223
rect -958 256913 298990 257223
rect -958 253913 298990 254223
rect -958 247913 298990 248223
rect -958 244913 298990 245223
rect -958 238913 298990 239223
rect -958 235913 298990 236223
rect -958 229913 298990 230223
rect -958 226913 298990 227223
rect -958 220913 298990 221223
rect -958 217913 298990 218223
rect -958 211913 298990 212223
rect -958 208913 298990 209223
rect -958 202913 298990 203223
rect -958 199913 298990 200223
rect -958 193913 298990 194223
rect -958 190913 298990 191223
rect -958 184913 298990 185223
rect -958 181913 298990 182223
rect -958 175913 298990 176223
rect -958 172913 298990 173223
rect -958 166913 298990 167223
rect -958 163913 298990 164223
rect -958 157913 298990 158223
rect -958 154913 298990 155223
rect -958 148913 298990 149223
rect -958 145913 298990 146223
rect -958 139913 298990 140223
rect -958 136913 298990 137223
rect -958 130913 298990 131223
rect -958 127913 298990 128223
rect -958 121913 298990 122223
rect -958 118913 298990 119223
rect -958 112913 298990 113223
rect -958 109913 298990 110223
rect -958 103913 298990 104223
rect -958 100913 298990 101223
rect -958 94913 298990 95223
rect -958 91913 298990 92223
rect -958 85913 298990 86223
rect -958 82913 298990 83223
rect -958 76913 298990 77223
rect -958 73913 298990 74223
rect -958 67913 298990 68223
rect -958 64913 298990 65223
rect -958 58913 298990 59223
rect -958 55913 298990 56223
rect -958 49913 298990 50223
rect -958 46913 298990 47223
rect -958 40913 298990 41223
rect -958 37913 298990 38223
rect -958 31913 298990 32223
rect -958 28913 298990 29223
rect -958 22913 298990 23223
rect -958 19913 298990 20223
rect -958 13913 298990 14223
rect -958 10913 298990 11223
rect -958 4913 298990 5223
rect -958 1913 298990 2223
rect -478 -342 298510 -32
rect -958 -822 298990 -512
<< labels >>
rlabel metal3 s 297780 120932 298500 121044 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal2 s 227164 297780 227276 298500 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 194236 297780 194348 298500 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 161308 297780 161420 298500 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 128380 297780 128492 298500 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 95452 297780 95564 298500 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 62524 297780 62636 298500 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 29596 297780 29708 298500 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal3 s -480 294364 240 294476 4 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s -480 272412 240 272524 4 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal3 s -480 250460 240 250572 4 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 297780 143332 298500 143444 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s -480 228508 240 228620 4 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s -480 206556 240 206668 4 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s -480 184604 240 184716 4 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal3 s -480 162652 240 162764 4 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s -480 140700 240 140812 4 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s -480 118748 240 118860 4 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s -480 96796 240 96908 4 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s -480 74844 240 74956 4 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s -480 52892 240 53004 4 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 297780 165732 298500 165844 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 297780 188132 298500 188244 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal3 s 297780 210532 298500 210644 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 297780 232932 298500 233044 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal3 s 297780 255332 298500 255444 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal3 s 297780 277732 298500 277844 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 293020 297780 293132 298500 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal2 s 260092 297780 260204 298500 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal3 s 297780 3332 298500 3444 6 io_in[0]
port 30 nsew signal input
rlabel metal3 s 297780 193732 298500 193844 6 io_in[10]
port 31 nsew signal input
rlabel metal3 s 297780 216132 298500 216244 6 io_in[11]
port 32 nsew signal input
rlabel metal3 s 297780 238532 298500 238644 6 io_in[12]
port 33 nsew signal input
rlabel metal3 s 297780 260932 298500 261044 6 io_in[13]
port 34 nsew signal input
rlabel metal3 s 297780 283332 298500 283444 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 284788 297780 284900 298500 6 io_in[15]
port 36 nsew signal input
rlabel metal2 s 251860 297780 251972 298500 6 io_in[16]
port 37 nsew signal input
rlabel metal2 s 218932 297780 219044 298500 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 186004 297780 186116 298500 6 io_in[18]
port 39 nsew signal input
rlabel metal2 s 153076 297780 153188 298500 6 io_in[19]
port 40 nsew signal input
rlabel metal3 s 297780 20132 298500 20244 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 120148 297780 120260 298500 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 87220 297780 87332 298500 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 54292 297780 54404 298500 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 21364 297780 21476 298500 6 io_in[23]
port 45 nsew signal input
rlabel metal3 s -480 288876 240 288988 4 io_in[24]
port 46 nsew signal input
rlabel metal3 s -480 266924 240 267036 4 io_in[25]
port 47 nsew signal input
rlabel metal3 s -480 244972 240 245084 4 io_in[26]
port 48 nsew signal input
rlabel metal3 s -480 223020 240 223132 4 io_in[27]
port 49 nsew signal input
rlabel metal3 s -480 201068 240 201180 4 io_in[28]
port 50 nsew signal input
rlabel metal3 s -480 179116 240 179228 4 io_in[29]
port 51 nsew signal input
rlabel metal3 s 297780 36932 298500 37044 6 io_in[2]
port 52 nsew signal input
rlabel metal3 s -480 157164 240 157276 4 io_in[30]
port 53 nsew signal input
rlabel metal3 s -480 135212 240 135324 4 io_in[31]
port 54 nsew signal input
rlabel metal3 s -480 113260 240 113372 4 io_in[32]
port 55 nsew signal input
rlabel metal3 s -480 91308 240 91420 4 io_in[33]
port 56 nsew signal input
rlabel metal3 s -480 69356 240 69468 4 io_in[34]
port 57 nsew signal input
rlabel metal3 s -480 47404 240 47516 4 io_in[35]
port 58 nsew signal input
rlabel metal3 s -480 30940 240 31052 4 io_in[36]
port 59 nsew signal input
rlabel metal3 s -480 14476 240 14588 4 io_in[37]
port 60 nsew signal input
rlabel metal3 s 297780 53732 298500 53844 6 io_in[3]
port 61 nsew signal input
rlabel metal3 s 297780 70532 298500 70644 6 io_in[4]
port 62 nsew signal input
rlabel metal3 s 297780 87332 298500 87444 6 io_in[5]
port 63 nsew signal input
rlabel metal3 s 297780 104132 298500 104244 6 io_in[6]
port 64 nsew signal input
rlabel metal3 s 297780 126532 298500 126644 6 io_in[7]
port 65 nsew signal input
rlabel metal3 s 297780 148932 298500 149044 6 io_in[8]
port 66 nsew signal input
rlabel metal3 s 297780 171332 298500 171444 6 io_in[9]
port 67 nsew signal input
rlabel metal3 s 297780 14532 298500 14644 6 io_oeb[0]
port 68 nsew signal output
rlabel metal3 s 297780 204932 298500 205044 6 io_oeb[10]
port 69 nsew signal output
rlabel metal3 s 297780 227332 298500 227444 6 io_oeb[11]
port 70 nsew signal output
rlabel metal3 s 297780 249732 298500 249844 6 io_oeb[12]
port 71 nsew signal output
rlabel metal3 s 297780 272132 298500 272244 6 io_oeb[13]
port 72 nsew signal output
rlabel metal3 s 297780 294532 298500 294644 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 268324 297780 268436 298500 6 io_oeb[15]
port 74 nsew signal output
rlabel metal2 s 235396 297780 235508 298500 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 202468 297780 202580 298500 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 169540 297780 169652 298500 6 io_oeb[18]
port 77 nsew signal output
rlabel metal2 s 136612 297780 136724 298500 6 io_oeb[19]
port 78 nsew signal output
rlabel metal3 s 297780 31332 298500 31444 6 io_oeb[1]
port 79 nsew signal output
rlabel metal2 s 103684 297780 103796 298500 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 70756 297780 70868 298500 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 37828 297780 37940 298500 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 4900 297780 5012 298500 6 io_oeb[23]
port 83 nsew signal output
rlabel metal3 s -480 277900 240 278012 4 io_oeb[24]
port 84 nsew signal output
rlabel metal3 s -480 255948 240 256060 4 io_oeb[25]
port 85 nsew signal output
rlabel metal3 s -480 233996 240 234108 4 io_oeb[26]
port 86 nsew signal output
rlabel metal3 s -480 212044 240 212156 4 io_oeb[27]
port 87 nsew signal output
rlabel metal3 s -480 190092 240 190204 4 io_oeb[28]
port 88 nsew signal output
rlabel metal3 s -480 168140 240 168252 4 io_oeb[29]
port 89 nsew signal output
rlabel metal3 s 297780 48132 298500 48244 6 io_oeb[2]
port 90 nsew signal output
rlabel metal3 s -480 146188 240 146300 4 io_oeb[30]
port 91 nsew signal output
rlabel metal3 s -480 124236 240 124348 4 io_oeb[31]
port 92 nsew signal output
rlabel metal3 s -480 102284 240 102396 4 io_oeb[32]
port 93 nsew signal output
rlabel metal3 s -480 80332 240 80444 4 io_oeb[33]
port 94 nsew signal output
rlabel metal3 s -480 58380 240 58492 4 io_oeb[34]
port 95 nsew signal output
rlabel metal3 s -480 36428 240 36540 4 io_oeb[35]
port 96 nsew signal output
rlabel metal3 s -480 19964 240 20076 4 io_oeb[36]
port 97 nsew signal output
rlabel metal3 s -480 3500 240 3612 4 io_oeb[37]
port 98 nsew signal output
rlabel metal3 s 297780 64932 298500 65044 6 io_oeb[3]
port 99 nsew signal output
rlabel metal3 s 297780 81732 298500 81844 6 io_oeb[4]
port 100 nsew signal output
rlabel metal3 s 297780 98532 298500 98644 6 io_oeb[5]
port 101 nsew signal output
rlabel metal3 s 297780 115332 298500 115444 6 io_oeb[6]
port 102 nsew signal output
rlabel metal3 s 297780 137732 298500 137844 6 io_oeb[7]
port 103 nsew signal output
rlabel metal3 s 297780 160132 298500 160244 6 io_oeb[8]
port 104 nsew signal output
rlabel metal3 s 297780 182532 298500 182644 6 io_oeb[9]
port 105 nsew signal output
rlabel metal3 s 297780 8932 298500 9044 6 io_out[0]
port 106 nsew signal output
rlabel metal3 s 297780 199332 298500 199444 6 io_out[10]
port 107 nsew signal output
rlabel metal3 s 297780 221732 298500 221844 6 io_out[11]
port 108 nsew signal output
rlabel metal3 s 297780 244132 298500 244244 6 io_out[12]
port 109 nsew signal output
rlabel metal3 s 297780 266532 298500 266644 6 io_out[13]
port 110 nsew signal output
rlabel metal3 s 297780 288932 298500 289044 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 276556 297780 276668 298500 6 io_out[15]
port 112 nsew signal output
rlabel metal2 s 243628 297780 243740 298500 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 210700 297780 210812 298500 6 io_out[17]
port 114 nsew signal output
rlabel metal2 s 177772 297780 177884 298500 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 144844 297780 144956 298500 6 io_out[19]
port 116 nsew signal output
rlabel metal3 s 297780 25732 298500 25844 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 111916 297780 112028 298500 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 78988 297780 79100 298500 6 io_out[21]
port 119 nsew signal output
rlabel metal2 s 46060 297780 46172 298500 6 io_out[22]
port 120 nsew signal output
rlabel metal2 s 13132 297780 13244 298500 6 io_out[23]
port 121 nsew signal output
rlabel metal3 s -480 283388 240 283500 4 io_out[24]
port 122 nsew signal output
rlabel metal3 s -480 261436 240 261548 4 io_out[25]
port 123 nsew signal output
rlabel metal3 s -480 239484 240 239596 4 io_out[26]
port 124 nsew signal output
rlabel metal3 s -480 217532 240 217644 4 io_out[27]
port 125 nsew signal output
rlabel metal3 s -480 195580 240 195692 4 io_out[28]
port 126 nsew signal output
rlabel metal3 s -480 173628 240 173740 4 io_out[29]
port 127 nsew signal output
rlabel metal3 s 297780 42532 298500 42644 6 io_out[2]
port 128 nsew signal output
rlabel metal3 s -480 151676 240 151788 4 io_out[30]
port 129 nsew signal output
rlabel metal3 s -480 129724 240 129836 4 io_out[31]
port 130 nsew signal output
rlabel metal3 s -480 107772 240 107884 4 io_out[32]
port 131 nsew signal output
rlabel metal3 s -480 85820 240 85932 4 io_out[33]
port 132 nsew signal output
rlabel metal3 s -480 63868 240 63980 4 io_out[34]
port 133 nsew signal output
rlabel metal3 s -480 41916 240 42028 4 io_out[35]
port 134 nsew signal output
rlabel metal3 s -480 25452 240 25564 4 io_out[36]
port 135 nsew signal output
rlabel metal3 s -480 8988 240 9100 4 io_out[37]
port 136 nsew signal output
rlabel metal3 s 297780 59332 298500 59444 6 io_out[3]
port 137 nsew signal output
rlabel metal3 s 297780 76132 298500 76244 6 io_out[4]
port 138 nsew signal output
rlabel metal3 s 297780 92932 298500 93044 6 io_out[5]
port 139 nsew signal output
rlabel metal3 s 297780 109732 298500 109844 6 io_out[6]
port 140 nsew signal output
rlabel metal3 s 297780 132132 298500 132244 6 io_out[7]
port 141 nsew signal output
rlabel metal3 s 297780 154532 298500 154644 6 io_out[8]
port 142 nsew signal output
rlabel metal3 s 297780 176932 298500 177044 6 io_out[9]
port 143 nsew signal output
rlabel metal2 s 70252 -480 70364 240 8 la_data_in[0]
port 144 nsew signal input
rlabel metal2 s 238252 -480 238364 240 8 la_data_in[100]
port 145 nsew signal input
rlabel metal2 s 239932 -480 240044 240 8 la_data_in[101]
port 146 nsew signal input
rlabel metal2 s 241612 -480 241724 240 8 la_data_in[102]
port 147 nsew signal input
rlabel metal2 s 243292 -480 243404 240 8 la_data_in[103]
port 148 nsew signal input
rlabel metal2 s 244972 -480 245084 240 8 la_data_in[104]
port 149 nsew signal input
rlabel metal2 s 246652 -480 246764 240 8 la_data_in[105]
port 150 nsew signal input
rlabel metal2 s 248332 -480 248444 240 8 la_data_in[106]
port 151 nsew signal input
rlabel metal2 s 250012 -480 250124 240 8 la_data_in[107]
port 152 nsew signal input
rlabel metal2 s 251692 -480 251804 240 8 la_data_in[108]
port 153 nsew signal input
rlabel metal2 s 253372 -480 253484 240 8 la_data_in[109]
port 154 nsew signal input
rlabel metal2 s 87052 -480 87164 240 8 la_data_in[10]
port 155 nsew signal input
rlabel metal2 s 255052 -480 255164 240 8 la_data_in[110]
port 156 nsew signal input
rlabel metal2 s 256732 -480 256844 240 8 la_data_in[111]
port 157 nsew signal input
rlabel metal2 s 258412 -480 258524 240 8 la_data_in[112]
port 158 nsew signal input
rlabel metal2 s 260092 -480 260204 240 8 la_data_in[113]
port 159 nsew signal input
rlabel metal2 s 261772 -480 261884 240 8 la_data_in[114]
port 160 nsew signal input
rlabel metal2 s 263452 -480 263564 240 8 la_data_in[115]
port 161 nsew signal input
rlabel metal2 s 265132 -480 265244 240 8 la_data_in[116]
port 162 nsew signal input
rlabel metal2 s 266812 -480 266924 240 8 la_data_in[117]
port 163 nsew signal input
rlabel metal2 s 268492 -480 268604 240 8 la_data_in[118]
port 164 nsew signal input
rlabel metal2 s 270172 -480 270284 240 8 la_data_in[119]
port 165 nsew signal input
rlabel metal2 s 88732 -480 88844 240 8 la_data_in[11]
port 166 nsew signal input
rlabel metal2 s 271852 -480 271964 240 8 la_data_in[120]
port 167 nsew signal input
rlabel metal2 s 273532 -480 273644 240 8 la_data_in[121]
port 168 nsew signal input
rlabel metal2 s 275212 -480 275324 240 8 la_data_in[122]
port 169 nsew signal input
rlabel metal2 s 276892 -480 277004 240 8 la_data_in[123]
port 170 nsew signal input
rlabel metal2 s 278572 -480 278684 240 8 la_data_in[124]
port 171 nsew signal input
rlabel metal2 s 280252 -480 280364 240 8 la_data_in[125]
port 172 nsew signal input
rlabel metal2 s 281932 -480 282044 240 8 la_data_in[126]
port 173 nsew signal input
rlabel metal2 s 283612 -480 283724 240 8 la_data_in[127]
port 174 nsew signal input
rlabel metal2 s 90412 -480 90524 240 8 la_data_in[12]
port 175 nsew signal input
rlabel metal2 s 92092 -480 92204 240 8 la_data_in[13]
port 176 nsew signal input
rlabel metal2 s 93772 -480 93884 240 8 la_data_in[14]
port 177 nsew signal input
rlabel metal2 s 95452 -480 95564 240 8 la_data_in[15]
port 178 nsew signal input
rlabel metal2 s 97132 -480 97244 240 8 la_data_in[16]
port 179 nsew signal input
rlabel metal2 s 98812 -480 98924 240 8 la_data_in[17]
port 180 nsew signal input
rlabel metal2 s 100492 -480 100604 240 8 la_data_in[18]
port 181 nsew signal input
rlabel metal2 s 102172 -480 102284 240 8 la_data_in[19]
port 182 nsew signal input
rlabel metal2 s 71932 -480 72044 240 8 la_data_in[1]
port 183 nsew signal input
rlabel metal2 s 103852 -480 103964 240 8 la_data_in[20]
port 184 nsew signal input
rlabel metal2 s 105532 -480 105644 240 8 la_data_in[21]
port 185 nsew signal input
rlabel metal2 s 107212 -480 107324 240 8 la_data_in[22]
port 186 nsew signal input
rlabel metal2 s 108892 -480 109004 240 8 la_data_in[23]
port 187 nsew signal input
rlabel metal2 s 110572 -480 110684 240 8 la_data_in[24]
port 188 nsew signal input
rlabel metal2 s 112252 -480 112364 240 8 la_data_in[25]
port 189 nsew signal input
rlabel metal2 s 113932 -480 114044 240 8 la_data_in[26]
port 190 nsew signal input
rlabel metal2 s 115612 -480 115724 240 8 la_data_in[27]
port 191 nsew signal input
rlabel metal2 s 117292 -480 117404 240 8 la_data_in[28]
port 192 nsew signal input
rlabel metal2 s 118972 -480 119084 240 8 la_data_in[29]
port 193 nsew signal input
rlabel metal2 s 73612 -480 73724 240 8 la_data_in[2]
port 194 nsew signal input
rlabel metal2 s 120652 -480 120764 240 8 la_data_in[30]
port 195 nsew signal input
rlabel metal2 s 122332 -480 122444 240 8 la_data_in[31]
port 196 nsew signal input
rlabel metal2 s 124012 -480 124124 240 8 la_data_in[32]
port 197 nsew signal input
rlabel metal2 s 125692 -480 125804 240 8 la_data_in[33]
port 198 nsew signal input
rlabel metal2 s 127372 -480 127484 240 8 la_data_in[34]
port 199 nsew signal input
rlabel metal2 s 129052 -480 129164 240 8 la_data_in[35]
port 200 nsew signal input
rlabel metal2 s 130732 -480 130844 240 8 la_data_in[36]
port 201 nsew signal input
rlabel metal2 s 132412 -480 132524 240 8 la_data_in[37]
port 202 nsew signal input
rlabel metal2 s 134092 -480 134204 240 8 la_data_in[38]
port 203 nsew signal input
rlabel metal2 s 135772 -480 135884 240 8 la_data_in[39]
port 204 nsew signal input
rlabel metal2 s 75292 -480 75404 240 8 la_data_in[3]
port 205 nsew signal input
rlabel metal2 s 137452 -480 137564 240 8 la_data_in[40]
port 206 nsew signal input
rlabel metal2 s 139132 -480 139244 240 8 la_data_in[41]
port 207 nsew signal input
rlabel metal2 s 140812 -480 140924 240 8 la_data_in[42]
port 208 nsew signal input
rlabel metal2 s 142492 -480 142604 240 8 la_data_in[43]
port 209 nsew signal input
rlabel metal2 s 144172 -480 144284 240 8 la_data_in[44]
port 210 nsew signal input
rlabel metal2 s 145852 -480 145964 240 8 la_data_in[45]
port 211 nsew signal input
rlabel metal2 s 147532 -480 147644 240 8 la_data_in[46]
port 212 nsew signal input
rlabel metal2 s 149212 -480 149324 240 8 la_data_in[47]
port 213 nsew signal input
rlabel metal2 s 150892 -480 151004 240 8 la_data_in[48]
port 214 nsew signal input
rlabel metal2 s 152572 -480 152684 240 8 la_data_in[49]
port 215 nsew signal input
rlabel metal2 s 76972 -480 77084 240 8 la_data_in[4]
port 216 nsew signal input
rlabel metal2 s 154252 -480 154364 240 8 la_data_in[50]
port 217 nsew signal input
rlabel metal2 s 155932 -480 156044 240 8 la_data_in[51]
port 218 nsew signal input
rlabel metal2 s 157612 -480 157724 240 8 la_data_in[52]
port 219 nsew signal input
rlabel metal2 s 159292 -480 159404 240 8 la_data_in[53]
port 220 nsew signal input
rlabel metal2 s 160972 -480 161084 240 8 la_data_in[54]
port 221 nsew signal input
rlabel metal2 s 162652 -480 162764 240 8 la_data_in[55]
port 222 nsew signal input
rlabel metal2 s 164332 -480 164444 240 8 la_data_in[56]
port 223 nsew signal input
rlabel metal2 s 166012 -480 166124 240 8 la_data_in[57]
port 224 nsew signal input
rlabel metal2 s 167692 -480 167804 240 8 la_data_in[58]
port 225 nsew signal input
rlabel metal2 s 169372 -480 169484 240 8 la_data_in[59]
port 226 nsew signal input
rlabel metal2 s 78652 -480 78764 240 8 la_data_in[5]
port 227 nsew signal input
rlabel metal2 s 171052 -480 171164 240 8 la_data_in[60]
port 228 nsew signal input
rlabel metal2 s 172732 -480 172844 240 8 la_data_in[61]
port 229 nsew signal input
rlabel metal2 s 174412 -480 174524 240 8 la_data_in[62]
port 230 nsew signal input
rlabel metal2 s 176092 -480 176204 240 8 la_data_in[63]
port 231 nsew signal input
rlabel metal2 s 177772 -480 177884 240 8 la_data_in[64]
port 232 nsew signal input
rlabel metal2 s 179452 -480 179564 240 8 la_data_in[65]
port 233 nsew signal input
rlabel metal2 s 181132 -480 181244 240 8 la_data_in[66]
port 234 nsew signal input
rlabel metal2 s 182812 -480 182924 240 8 la_data_in[67]
port 235 nsew signal input
rlabel metal2 s 184492 -480 184604 240 8 la_data_in[68]
port 236 nsew signal input
rlabel metal2 s 186172 -480 186284 240 8 la_data_in[69]
port 237 nsew signal input
rlabel metal2 s 80332 -480 80444 240 8 la_data_in[6]
port 238 nsew signal input
rlabel metal2 s 187852 -480 187964 240 8 la_data_in[70]
port 239 nsew signal input
rlabel metal2 s 189532 -480 189644 240 8 la_data_in[71]
port 240 nsew signal input
rlabel metal2 s 191212 -480 191324 240 8 la_data_in[72]
port 241 nsew signal input
rlabel metal2 s 192892 -480 193004 240 8 la_data_in[73]
port 242 nsew signal input
rlabel metal2 s 194572 -480 194684 240 8 la_data_in[74]
port 243 nsew signal input
rlabel metal2 s 196252 -480 196364 240 8 la_data_in[75]
port 244 nsew signal input
rlabel metal2 s 197932 -480 198044 240 8 la_data_in[76]
port 245 nsew signal input
rlabel metal2 s 199612 -480 199724 240 8 la_data_in[77]
port 246 nsew signal input
rlabel metal2 s 201292 -480 201404 240 8 la_data_in[78]
port 247 nsew signal input
rlabel metal2 s 202972 -480 203084 240 8 la_data_in[79]
port 248 nsew signal input
rlabel metal2 s 82012 -480 82124 240 8 la_data_in[7]
port 249 nsew signal input
rlabel metal2 s 204652 -480 204764 240 8 la_data_in[80]
port 250 nsew signal input
rlabel metal2 s 206332 -480 206444 240 8 la_data_in[81]
port 251 nsew signal input
rlabel metal2 s 208012 -480 208124 240 8 la_data_in[82]
port 252 nsew signal input
rlabel metal2 s 209692 -480 209804 240 8 la_data_in[83]
port 253 nsew signal input
rlabel metal2 s 211372 -480 211484 240 8 la_data_in[84]
port 254 nsew signal input
rlabel metal2 s 213052 -480 213164 240 8 la_data_in[85]
port 255 nsew signal input
rlabel metal2 s 214732 -480 214844 240 8 la_data_in[86]
port 256 nsew signal input
rlabel metal2 s 216412 -480 216524 240 8 la_data_in[87]
port 257 nsew signal input
rlabel metal2 s 218092 -480 218204 240 8 la_data_in[88]
port 258 nsew signal input
rlabel metal2 s 219772 -480 219884 240 8 la_data_in[89]
port 259 nsew signal input
rlabel metal2 s 83692 -480 83804 240 8 la_data_in[8]
port 260 nsew signal input
rlabel metal2 s 221452 -480 221564 240 8 la_data_in[90]
port 261 nsew signal input
rlabel metal2 s 223132 -480 223244 240 8 la_data_in[91]
port 262 nsew signal input
rlabel metal2 s 224812 -480 224924 240 8 la_data_in[92]
port 263 nsew signal input
rlabel metal2 s 226492 -480 226604 240 8 la_data_in[93]
port 264 nsew signal input
rlabel metal2 s 228172 -480 228284 240 8 la_data_in[94]
port 265 nsew signal input
rlabel metal2 s 229852 -480 229964 240 8 la_data_in[95]
port 266 nsew signal input
rlabel metal2 s 231532 -480 231644 240 8 la_data_in[96]
port 267 nsew signal input
rlabel metal2 s 233212 -480 233324 240 8 la_data_in[97]
port 268 nsew signal input
rlabel metal2 s 234892 -480 235004 240 8 la_data_in[98]
port 269 nsew signal input
rlabel metal2 s 236572 -480 236684 240 8 la_data_in[99]
port 270 nsew signal input
rlabel metal2 s 85372 -480 85484 240 8 la_data_in[9]
port 271 nsew signal input
rlabel metal2 s 70812 -480 70924 240 8 la_data_out[0]
port 272 nsew signal output
rlabel metal2 s 238812 -480 238924 240 8 la_data_out[100]
port 273 nsew signal output
rlabel metal2 s 240492 -480 240604 240 8 la_data_out[101]
port 274 nsew signal output
rlabel metal2 s 242172 -480 242284 240 8 la_data_out[102]
port 275 nsew signal output
rlabel metal2 s 243852 -480 243964 240 8 la_data_out[103]
port 276 nsew signal output
rlabel metal2 s 245532 -480 245644 240 8 la_data_out[104]
port 277 nsew signal output
rlabel metal2 s 247212 -480 247324 240 8 la_data_out[105]
port 278 nsew signal output
rlabel metal2 s 248892 -480 249004 240 8 la_data_out[106]
port 279 nsew signal output
rlabel metal2 s 250572 -480 250684 240 8 la_data_out[107]
port 280 nsew signal output
rlabel metal2 s 252252 -480 252364 240 8 la_data_out[108]
port 281 nsew signal output
rlabel metal2 s 253932 -480 254044 240 8 la_data_out[109]
port 282 nsew signal output
rlabel metal2 s 87612 -480 87724 240 8 la_data_out[10]
port 283 nsew signal output
rlabel metal2 s 255612 -480 255724 240 8 la_data_out[110]
port 284 nsew signal output
rlabel metal2 s 257292 -480 257404 240 8 la_data_out[111]
port 285 nsew signal output
rlabel metal2 s 258972 -480 259084 240 8 la_data_out[112]
port 286 nsew signal output
rlabel metal2 s 260652 -480 260764 240 8 la_data_out[113]
port 287 nsew signal output
rlabel metal2 s 262332 -480 262444 240 8 la_data_out[114]
port 288 nsew signal output
rlabel metal2 s 264012 -480 264124 240 8 la_data_out[115]
port 289 nsew signal output
rlabel metal2 s 265692 -480 265804 240 8 la_data_out[116]
port 290 nsew signal output
rlabel metal2 s 267372 -480 267484 240 8 la_data_out[117]
port 291 nsew signal output
rlabel metal2 s 269052 -480 269164 240 8 la_data_out[118]
port 292 nsew signal output
rlabel metal2 s 270732 -480 270844 240 8 la_data_out[119]
port 293 nsew signal output
rlabel metal2 s 89292 -480 89404 240 8 la_data_out[11]
port 294 nsew signal output
rlabel metal2 s 272412 -480 272524 240 8 la_data_out[120]
port 295 nsew signal output
rlabel metal2 s 274092 -480 274204 240 8 la_data_out[121]
port 296 nsew signal output
rlabel metal2 s 275772 -480 275884 240 8 la_data_out[122]
port 297 nsew signal output
rlabel metal2 s 277452 -480 277564 240 8 la_data_out[123]
port 298 nsew signal output
rlabel metal2 s 279132 -480 279244 240 8 la_data_out[124]
port 299 nsew signal output
rlabel metal2 s 280812 -480 280924 240 8 la_data_out[125]
port 300 nsew signal output
rlabel metal2 s 282492 -480 282604 240 8 la_data_out[126]
port 301 nsew signal output
rlabel metal2 s 284172 -480 284284 240 8 la_data_out[127]
port 302 nsew signal output
rlabel metal2 s 90972 -480 91084 240 8 la_data_out[12]
port 303 nsew signal output
rlabel metal2 s 92652 -480 92764 240 8 la_data_out[13]
port 304 nsew signal output
rlabel metal2 s 94332 -480 94444 240 8 la_data_out[14]
port 305 nsew signal output
rlabel metal2 s 96012 -480 96124 240 8 la_data_out[15]
port 306 nsew signal output
rlabel metal2 s 97692 -480 97804 240 8 la_data_out[16]
port 307 nsew signal output
rlabel metal2 s 99372 -480 99484 240 8 la_data_out[17]
port 308 nsew signal output
rlabel metal2 s 101052 -480 101164 240 8 la_data_out[18]
port 309 nsew signal output
rlabel metal2 s 102732 -480 102844 240 8 la_data_out[19]
port 310 nsew signal output
rlabel metal2 s 72492 -480 72604 240 8 la_data_out[1]
port 311 nsew signal output
rlabel metal2 s 104412 -480 104524 240 8 la_data_out[20]
port 312 nsew signal output
rlabel metal2 s 106092 -480 106204 240 8 la_data_out[21]
port 313 nsew signal output
rlabel metal2 s 107772 -480 107884 240 8 la_data_out[22]
port 314 nsew signal output
rlabel metal2 s 109452 -480 109564 240 8 la_data_out[23]
port 315 nsew signal output
rlabel metal2 s 111132 -480 111244 240 8 la_data_out[24]
port 316 nsew signal output
rlabel metal2 s 112812 -480 112924 240 8 la_data_out[25]
port 317 nsew signal output
rlabel metal2 s 114492 -480 114604 240 8 la_data_out[26]
port 318 nsew signal output
rlabel metal2 s 116172 -480 116284 240 8 la_data_out[27]
port 319 nsew signal output
rlabel metal2 s 117852 -480 117964 240 8 la_data_out[28]
port 320 nsew signal output
rlabel metal2 s 119532 -480 119644 240 8 la_data_out[29]
port 321 nsew signal output
rlabel metal2 s 74172 -480 74284 240 8 la_data_out[2]
port 322 nsew signal output
rlabel metal2 s 121212 -480 121324 240 8 la_data_out[30]
port 323 nsew signal output
rlabel metal2 s 122892 -480 123004 240 8 la_data_out[31]
port 324 nsew signal output
rlabel metal2 s 124572 -480 124684 240 8 la_data_out[32]
port 325 nsew signal output
rlabel metal2 s 126252 -480 126364 240 8 la_data_out[33]
port 326 nsew signal output
rlabel metal2 s 127932 -480 128044 240 8 la_data_out[34]
port 327 nsew signal output
rlabel metal2 s 129612 -480 129724 240 8 la_data_out[35]
port 328 nsew signal output
rlabel metal2 s 131292 -480 131404 240 8 la_data_out[36]
port 329 nsew signal output
rlabel metal2 s 132972 -480 133084 240 8 la_data_out[37]
port 330 nsew signal output
rlabel metal2 s 134652 -480 134764 240 8 la_data_out[38]
port 331 nsew signal output
rlabel metal2 s 136332 -480 136444 240 8 la_data_out[39]
port 332 nsew signal output
rlabel metal2 s 75852 -480 75964 240 8 la_data_out[3]
port 333 nsew signal output
rlabel metal2 s 138012 -480 138124 240 8 la_data_out[40]
port 334 nsew signal output
rlabel metal2 s 139692 -480 139804 240 8 la_data_out[41]
port 335 nsew signal output
rlabel metal2 s 141372 -480 141484 240 8 la_data_out[42]
port 336 nsew signal output
rlabel metal2 s 143052 -480 143164 240 8 la_data_out[43]
port 337 nsew signal output
rlabel metal2 s 144732 -480 144844 240 8 la_data_out[44]
port 338 nsew signal output
rlabel metal2 s 146412 -480 146524 240 8 la_data_out[45]
port 339 nsew signal output
rlabel metal2 s 148092 -480 148204 240 8 la_data_out[46]
port 340 nsew signal output
rlabel metal2 s 149772 -480 149884 240 8 la_data_out[47]
port 341 nsew signal output
rlabel metal2 s 151452 -480 151564 240 8 la_data_out[48]
port 342 nsew signal output
rlabel metal2 s 153132 -480 153244 240 8 la_data_out[49]
port 343 nsew signal output
rlabel metal2 s 77532 -480 77644 240 8 la_data_out[4]
port 344 nsew signal output
rlabel metal2 s 154812 -480 154924 240 8 la_data_out[50]
port 345 nsew signal output
rlabel metal2 s 156492 -480 156604 240 8 la_data_out[51]
port 346 nsew signal output
rlabel metal2 s 158172 -480 158284 240 8 la_data_out[52]
port 347 nsew signal output
rlabel metal2 s 159852 -480 159964 240 8 la_data_out[53]
port 348 nsew signal output
rlabel metal2 s 161532 -480 161644 240 8 la_data_out[54]
port 349 nsew signal output
rlabel metal2 s 163212 -480 163324 240 8 la_data_out[55]
port 350 nsew signal output
rlabel metal2 s 164892 -480 165004 240 8 la_data_out[56]
port 351 nsew signal output
rlabel metal2 s 166572 -480 166684 240 8 la_data_out[57]
port 352 nsew signal output
rlabel metal2 s 168252 -480 168364 240 8 la_data_out[58]
port 353 nsew signal output
rlabel metal2 s 169932 -480 170044 240 8 la_data_out[59]
port 354 nsew signal output
rlabel metal2 s 79212 -480 79324 240 8 la_data_out[5]
port 355 nsew signal output
rlabel metal2 s 171612 -480 171724 240 8 la_data_out[60]
port 356 nsew signal output
rlabel metal2 s 173292 -480 173404 240 8 la_data_out[61]
port 357 nsew signal output
rlabel metal2 s 174972 -480 175084 240 8 la_data_out[62]
port 358 nsew signal output
rlabel metal2 s 176652 -480 176764 240 8 la_data_out[63]
port 359 nsew signal output
rlabel metal2 s 178332 -480 178444 240 8 la_data_out[64]
port 360 nsew signal output
rlabel metal2 s 180012 -480 180124 240 8 la_data_out[65]
port 361 nsew signal output
rlabel metal2 s 181692 -480 181804 240 8 la_data_out[66]
port 362 nsew signal output
rlabel metal2 s 183372 -480 183484 240 8 la_data_out[67]
port 363 nsew signal output
rlabel metal2 s 185052 -480 185164 240 8 la_data_out[68]
port 364 nsew signal output
rlabel metal2 s 186732 -480 186844 240 8 la_data_out[69]
port 365 nsew signal output
rlabel metal2 s 80892 -480 81004 240 8 la_data_out[6]
port 366 nsew signal output
rlabel metal2 s 188412 -480 188524 240 8 la_data_out[70]
port 367 nsew signal output
rlabel metal2 s 190092 -480 190204 240 8 la_data_out[71]
port 368 nsew signal output
rlabel metal2 s 191772 -480 191884 240 8 la_data_out[72]
port 369 nsew signal output
rlabel metal2 s 193452 -480 193564 240 8 la_data_out[73]
port 370 nsew signal output
rlabel metal2 s 195132 -480 195244 240 8 la_data_out[74]
port 371 nsew signal output
rlabel metal2 s 196812 -480 196924 240 8 la_data_out[75]
port 372 nsew signal output
rlabel metal2 s 198492 -480 198604 240 8 la_data_out[76]
port 373 nsew signal output
rlabel metal2 s 200172 -480 200284 240 8 la_data_out[77]
port 374 nsew signal output
rlabel metal2 s 201852 -480 201964 240 8 la_data_out[78]
port 375 nsew signal output
rlabel metal2 s 203532 -480 203644 240 8 la_data_out[79]
port 376 nsew signal output
rlabel metal2 s 82572 -480 82684 240 8 la_data_out[7]
port 377 nsew signal output
rlabel metal2 s 205212 -480 205324 240 8 la_data_out[80]
port 378 nsew signal output
rlabel metal2 s 206892 -480 207004 240 8 la_data_out[81]
port 379 nsew signal output
rlabel metal2 s 208572 -480 208684 240 8 la_data_out[82]
port 380 nsew signal output
rlabel metal2 s 210252 -480 210364 240 8 la_data_out[83]
port 381 nsew signal output
rlabel metal2 s 211932 -480 212044 240 8 la_data_out[84]
port 382 nsew signal output
rlabel metal2 s 213612 -480 213724 240 8 la_data_out[85]
port 383 nsew signal output
rlabel metal2 s 215292 -480 215404 240 8 la_data_out[86]
port 384 nsew signal output
rlabel metal2 s 216972 -480 217084 240 8 la_data_out[87]
port 385 nsew signal output
rlabel metal2 s 218652 -480 218764 240 8 la_data_out[88]
port 386 nsew signal output
rlabel metal2 s 220332 -480 220444 240 8 la_data_out[89]
port 387 nsew signal output
rlabel metal2 s 84252 -480 84364 240 8 la_data_out[8]
port 388 nsew signal output
rlabel metal2 s 222012 -480 222124 240 8 la_data_out[90]
port 389 nsew signal output
rlabel metal2 s 223692 -480 223804 240 8 la_data_out[91]
port 390 nsew signal output
rlabel metal2 s 225372 -480 225484 240 8 la_data_out[92]
port 391 nsew signal output
rlabel metal2 s 227052 -480 227164 240 8 la_data_out[93]
port 392 nsew signal output
rlabel metal2 s 228732 -480 228844 240 8 la_data_out[94]
port 393 nsew signal output
rlabel metal2 s 230412 -480 230524 240 8 la_data_out[95]
port 394 nsew signal output
rlabel metal2 s 232092 -480 232204 240 8 la_data_out[96]
port 395 nsew signal output
rlabel metal2 s 233772 -480 233884 240 8 la_data_out[97]
port 396 nsew signal output
rlabel metal2 s 235452 -480 235564 240 8 la_data_out[98]
port 397 nsew signal output
rlabel metal2 s 237132 -480 237244 240 8 la_data_out[99]
port 398 nsew signal output
rlabel metal2 s 85932 -480 86044 240 8 la_data_out[9]
port 399 nsew signal output
rlabel metal2 s 71372 -480 71484 240 8 la_oenb[0]
port 400 nsew signal input
rlabel metal2 s 239372 -480 239484 240 8 la_oenb[100]
port 401 nsew signal input
rlabel metal2 s 241052 -480 241164 240 8 la_oenb[101]
port 402 nsew signal input
rlabel metal2 s 242732 -480 242844 240 8 la_oenb[102]
port 403 nsew signal input
rlabel metal2 s 244412 -480 244524 240 8 la_oenb[103]
port 404 nsew signal input
rlabel metal2 s 246092 -480 246204 240 8 la_oenb[104]
port 405 nsew signal input
rlabel metal2 s 247772 -480 247884 240 8 la_oenb[105]
port 406 nsew signal input
rlabel metal2 s 249452 -480 249564 240 8 la_oenb[106]
port 407 nsew signal input
rlabel metal2 s 251132 -480 251244 240 8 la_oenb[107]
port 408 nsew signal input
rlabel metal2 s 252812 -480 252924 240 8 la_oenb[108]
port 409 nsew signal input
rlabel metal2 s 254492 -480 254604 240 8 la_oenb[109]
port 410 nsew signal input
rlabel metal2 s 88172 -480 88284 240 8 la_oenb[10]
port 411 nsew signal input
rlabel metal2 s 256172 -480 256284 240 8 la_oenb[110]
port 412 nsew signal input
rlabel metal2 s 257852 -480 257964 240 8 la_oenb[111]
port 413 nsew signal input
rlabel metal2 s 259532 -480 259644 240 8 la_oenb[112]
port 414 nsew signal input
rlabel metal2 s 261212 -480 261324 240 8 la_oenb[113]
port 415 nsew signal input
rlabel metal2 s 262892 -480 263004 240 8 la_oenb[114]
port 416 nsew signal input
rlabel metal2 s 264572 -480 264684 240 8 la_oenb[115]
port 417 nsew signal input
rlabel metal2 s 266252 -480 266364 240 8 la_oenb[116]
port 418 nsew signal input
rlabel metal2 s 267932 -480 268044 240 8 la_oenb[117]
port 419 nsew signal input
rlabel metal2 s 269612 -480 269724 240 8 la_oenb[118]
port 420 nsew signal input
rlabel metal2 s 271292 -480 271404 240 8 la_oenb[119]
port 421 nsew signal input
rlabel metal2 s 89852 -480 89964 240 8 la_oenb[11]
port 422 nsew signal input
rlabel metal2 s 272972 -480 273084 240 8 la_oenb[120]
port 423 nsew signal input
rlabel metal2 s 274652 -480 274764 240 8 la_oenb[121]
port 424 nsew signal input
rlabel metal2 s 276332 -480 276444 240 8 la_oenb[122]
port 425 nsew signal input
rlabel metal2 s 278012 -480 278124 240 8 la_oenb[123]
port 426 nsew signal input
rlabel metal2 s 279692 -480 279804 240 8 la_oenb[124]
port 427 nsew signal input
rlabel metal2 s 281372 -480 281484 240 8 la_oenb[125]
port 428 nsew signal input
rlabel metal2 s 283052 -480 283164 240 8 la_oenb[126]
port 429 nsew signal input
rlabel metal2 s 284732 -480 284844 240 8 la_oenb[127]
port 430 nsew signal input
rlabel metal2 s 91532 -480 91644 240 8 la_oenb[12]
port 431 nsew signal input
rlabel metal2 s 93212 -480 93324 240 8 la_oenb[13]
port 432 nsew signal input
rlabel metal2 s 94892 -480 95004 240 8 la_oenb[14]
port 433 nsew signal input
rlabel metal2 s 96572 -480 96684 240 8 la_oenb[15]
port 434 nsew signal input
rlabel metal2 s 98252 -480 98364 240 8 la_oenb[16]
port 435 nsew signal input
rlabel metal2 s 99932 -480 100044 240 8 la_oenb[17]
port 436 nsew signal input
rlabel metal2 s 101612 -480 101724 240 8 la_oenb[18]
port 437 nsew signal input
rlabel metal2 s 103292 -480 103404 240 8 la_oenb[19]
port 438 nsew signal input
rlabel metal2 s 73052 -480 73164 240 8 la_oenb[1]
port 439 nsew signal input
rlabel metal2 s 104972 -480 105084 240 8 la_oenb[20]
port 440 nsew signal input
rlabel metal2 s 106652 -480 106764 240 8 la_oenb[21]
port 441 nsew signal input
rlabel metal2 s 108332 -480 108444 240 8 la_oenb[22]
port 442 nsew signal input
rlabel metal2 s 110012 -480 110124 240 8 la_oenb[23]
port 443 nsew signal input
rlabel metal2 s 111692 -480 111804 240 8 la_oenb[24]
port 444 nsew signal input
rlabel metal2 s 113372 -480 113484 240 8 la_oenb[25]
port 445 nsew signal input
rlabel metal2 s 115052 -480 115164 240 8 la_oenb[26]
port 446 nsew signal input
rlabel metal2 s 116732 -480 116844 240 8 la_oenb[27]
port 447 nsew signal input
rlabel metal2 s 118412 -480 118524 240 8 la_oenb[28]
port 448 nsew signal input
rlabel metal2 s 120092 -480 120204 240 8 la_oenb[29]
port 449 nsew signal input
rlabel metal2 s 74732 -480 74844 240 8 la_oenb[2]
port 450 nsew signal input
rlabel metal2 s 121772 -480 121884 240 8 la_oenb[30]
port 451 nsew signal input
rlabel metal2 s 123452 -480 123564 240 8 la_oenb[31]
port 452 nsew signal input
rlabel metal2 s 125132 -480 125244 240 8 la_oenb[32]
port 453 nsew signal input
rlabel metal2 s 126812 -480 126924 240 8 la_oenb[33]
port 454 nsew signal input
rlabel metal2 s 128492 -480 128604 240 8 la_oenb[34]
port 455 nsew signal input
rlabel metal2 s 130172 -480 130284 240 8 la_oenb[35]
port 456 nsew signal input
rlabel metal2 s 131852 -480 131964 240 8 la_oenb[36]
port 457 nsew signal input
rlabel metal2 s 133532 -480 133644 240 8 la_oenb[37]
port 458 nsew signal input
rlabel metal2 s 135212 -480 135324 240 8 la_oenb[38]
port 459 nsew signal input
rlabel metal2 s 136892 -480 137004 240 8 la_oenb[39]
port 460 nsew signal input
rlabel metal2 s 76412 -480 76524 240 8 la_oenb[3]
port 461 nsew signal input
rlabel metal2 s 138572 -480 138684 240 8 la_oenb[40]
port 462 nsew signal input
rlabel metal2 s 140252 -480 140364 240 8 la_oenb[41]
port 463 nsew signal input
rlabel metal2 s 141932 -480 142044 240 8 la_oenb[42]
port 464 nsew signal input
rlabel metal2 s 143612 -480 143724 240 8 la_oenb[43]
port 465 nsew signal input
rlabel metal2 s 145292 -480 145404 240 8 la_oenb[44]
port 466 nsew signal input
rlabel metal2 s 146972 -480 147084 240 8 la_oenb[45]
port 467 nsew signal input
rlabel metal2 s 148652 -480 148764 240 8 la_oenb[46]
port 468 nsew signal input
rlabel metal2 s 150332 -480 150444 240 8 la_oenb[47]
port 469 nsew signal input
rlabel metal2 s 152012 -480 152124 240 8 la_oenb[48]
port 470 nsew signal input
rlabel metal2 s 153692 -480 153804 240 8 la_oenb[49]
port 471 nsew signal input
rlabel metal2 s 78092 -480 78204 240 8 la_oenb[4]
port 472 nsew signal input
rlabel metal2 s 155372 -480 155484 240 8 la_oenb[50]
port 473 nsew signal input
rlabel metal2 s 157052 -480 157164 240 8 la_oenb[51]
port 474 nsew signal input
rlabel metal2 s 158732 -480 158844 240 8 la_oenb[52]
port 475 nsew signal input
rlabel metal2 s 160412 -480 160524 240 8 la_oenb[53]
port 476 nsew signal input
rlabel metal2 s 162092 -480 162204 240 8 la_oenb[54]
port 477 nsew signal input
rlabel metal2 s 163772 -480 163884 240 8 la_oenb[55]
port 478 nsew signal input
rlabel metal2 s 165452 -480 165564 240 8 la_oenb[56]
port 479 nsew signal input
rlabel metal2 s 167132 -480 167244 240 8 la_oenb[57]
port 480 nsew signal input
rlabel metal2 s 168812 -480 168924 240 8 la_oenb[58]
port 481 nsew signal input
rlabel metal2 s 170492 -480 170604 240 8 la_oenb[59]
port 482 nsew signal input
rlabel metal2 s 79772 -480 79884 240 8 la_oenb[5]
port 483 nsew signal input
rlabel metal2 s 172172 -480 172284 240 8 la_oenb[60]
port 484 nsew signal input
rlabel metal2 s 173852 -480 173964 240 8 la_oenb[61]
port 485 nsew signal input
rlabel metal2 s 175532 -480 175644 240 8 la_oenb[62]
port 486 nsew signal input
rlabel metal2 s 177212 -480 177324 240 8 la_oenb[63]
port 487 nsew signal input
rlabel metal2 s 178892 -480 179004 240 8 la_oenb[64]
port 488 nsew signal input
rlabel metal2 s 180572 -480 180684 240 8 la_oenb[65]
port 489 nsew signal input
rlabel metal2 s 182252 -480 182364 240 8 la_oenb[66]
port 490 nsew signal input
rlabel metal2 s 183932 -480 184044 240 8 la_oenb[67]
port 491 nsew signal input
rlabel metal2 s 185612 -480 185724 240 8 la_oenb[68]
port 492 nsew signal input
rlabel metal2 s 187292 -480 187404 240 8 la_oenb[69]
port 493 nsew signal input
rlabel metal2 s 81452 -480 81564 240 8 la_oenb[6]
port 494 nsew signal input
rlabel metal2 s 188972 -480 189084 240 8 la_oenb[70]
port 495 nsew signal input
rlabel metal2 s 190652 -480 190764 240 8 la_oenb[71]
port 496 nsew signal input
rlabel metal2 s 192332 -480 192444 240 8 la_oenb[72]
port 497 nsew signal input
rlabel metal2 s 194012 -480 194124 240 8 la_oenb[73]
port 498 nsew signal input
rlabel metal2 s 195692 -480 195804 240 8 la_oenb[74]
port 499 nsew signal input
rlabel metal2 s 197372 -480 197484 240 8 la_oenb[75]
port 500 nsew signal input
rlabel metal2 s 199052 -480 199164 240 8 la_oenb[76]
port 501 nsew signal input
rlabel metal2 s 200732 -480 200844 240 8 la_oenb[77]
port 502 nsew signal input
rlabel metal2 s 202412 -480 202524 240 8 la_oenb[78]
port 503 nsew signal input
rlabel metal2 s 204092 -480 204204 240 8 la_oenb[79]
port 504 nsew signal input
rlabel metal2 s 83132 -480 83244 240 8 la_oenb[7]
port 505 nsew signal input
rlabel metal2 s 205772 -480 205884 240 8 la_oenb[80]
port 506 nsew signal input
rlabel metal2 s 207452 -480 207564 240 8 la_oenb[81]
port 507 nsew signal input
rlabel metal2 s 209132 -480 209244 240 8 la_oenb[82]
port 508 nsew signal input
rlabel metal2 s 210812 -480 210924 240 8 la_oenb[83]
port 509 nsew signal input
rlabel metal2 s 212492 -480 212604 240 8 la_oenb[84]
port 510 nsew signal input
rlabel metal2 s 214172 -480 214284 240 8 la_oenb[85]
port 511 nsew signal input
rlabel metal2 s 215852 -480 215964 240 8 la_oenb[86]
port 512 nsew signal input
rlabel metal2 s 217532 -480 217644 240 8 la_oenb[87]
port 513 nsew signal input
rlabel metal2 s 219212 -480 219324 240 8 la_oenb[88]
port 514 nsew signal input
rlabel metal2 s 220892 -480 221004 240 8 la_oenb[89]
port 515 nsew signal input
rlabel metal2 s 84812 -480 84924 240 8 la_oenb[8]
port 516 nsew signal input
rlabel metal2 s 222572 -480 222684 240 8 la_oenb[90]
port 517 nsew signal input
rlabel metal2 s 224252 -480 224364 240 8 la_oenb[91]
port 518 nsew signal input
rlabel metal2 s 225932 -480 226044 240 8 la_oenb[92]
port 519 nsew signal input
rlabel metal2 s 227612 -480 227724 240 8 la_oenb[93]
port 520 nsew signal input
rlabel metal2 s 229292 -480 229404 240 8 la_oenb[94]
port 521 nsew signal input
rlabel metal2 s 230972 -480 231084 240 8 la_oenb[95]
port 522 nsew signal input
rlabel metal2 s 232652 -480 232764 240 8 la_oenb[96]
port 523 nsew signal input
rlabel metal2 s 234332 -480 234444 240 8 la_oenb[97]
port 524 nsew signal input
rlabel metal2 s 236012 -480 236124 240 8 la_oenb[98]
port 525 nsew signal input
rlabel metal2 s 237692 -480 237804 240 8 la_oenb[99]
port 526 nsew signal input
rlabel metal2 s 86492 -480 86604 240 8 la_oenb[9]
port 527 nsew signal input
rlabel metal2 s 285292 -480 285404 240 8 user_clock2
port 528 nsew signal input
rlabel metal2 s 285852 -480 285964 240 8 user_irq[0]
port 529 nsew signal output
rlabel metal2 s 286412 -480 286524 240 8 user_irq[1]
port 530 nsew signal output
rlabel metal2 s 286972 -480 287084 240 8 user_irq[2]
port 531 nsew signal output
rlabel metal4 s -478 -342 -168 298654 4 vdd
port 532 nsew power bidirectional
rlabel metal5 s -478 -342 298510 -32 8 vdd
port 532 nsew power bidirectional
rlabel metal5 s -478 298344 298510 298654 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 298200 -342 298510 298654 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 1577 -822 1887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 10577 -822 10887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 19577 -822 19887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 28577 -822 28887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 37577 -822 37887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 46577 -822 46887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 55577 -822 55887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 64577 -822 64887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 73577 -822 73887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 82577 -822 82887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 91577 -822 91887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 100577 -822 100887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 109577 -822 109887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 118577 -822 118887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 127577 -822 127887 169510 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 127577 228466 127887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 136577 -822 136887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 145577 -822 145887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 154577 -822 154887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 163577 -822 163887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 172577 -822 172887 224765 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 172577 228091 172887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 181577 -822 181887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 190577 -822 190887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 199577 -822 199887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 208577 -822 208887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 217577 -822 217887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 226577 -822 226887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 235577 -822 235887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 244577 -822 244887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 253577 -822 253887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 262577 -822 262887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 271577 -822 271887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 280577 -822 280887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s 289577 -822 289887 299134 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 1913 298990 2223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 10913 298990 11223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 19913 298990 20223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 28913 298990 29223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 37913 298990 38223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 46913 298990 47223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 55913 298990 56223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 64913 298990 65223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 73913 298990 74223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 82913 298990 83223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 91913 298990 92223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 100913 298990 101223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 109913 298990 110223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 118913 298990 119223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 127913 298990 128223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 136913 298990 137223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 145913 298990 146223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 154913 298990 155223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 163913 298990 164223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 172913 298990 173223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 181913 298990 182223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 190913 298990 191223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 199913 298990 200223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 208913 298990 209223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 217913 298990 218223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 226913 298990 227223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 235913 298990 236223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 244913 298990 245223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 253913 298990 254223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 262913 298990 263223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 271913 298990 272223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 280913 298990 281223 6 vdd
port 532 nsew power bidirectional
rlabel metal5 s -958 289913 298990 290223 6 vdd
port 532 nsew power bidirectional
rlabel metal4 s -958 -822 -648 299134 4 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 -822 298990 -512 8 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 298824 298990 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 298680 -822 298990 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 3437 -822 3747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 12437 -822 12747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 21437 -822 21747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 30437 -822 30747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 39437 -822 39747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 48437 -822 48747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 57437 -822 57747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 66437 -822 66747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 75437 -822 75747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 84437 -822 84747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 93437 -822 93747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 102437 -822 102747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 111437 -822 111747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 120437 -822 120747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 129437 -822 129747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 138437 -822 138747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 147437 -822 147747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 156437 -822 156747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 165437 -822 165747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 174437 -822 174747 224765 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 174437 228091 174747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 183437 -822 183747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 192437 -822 192747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 201437 -822 201747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 210437 -822 210747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 219437 -822 219747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 228437 -822 228747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 237437 -822 237747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 246437 -822 246747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 255437 -822 255747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 264437 -822 264747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 273437 -822 273747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 282437 -822 282747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal4 s 291437 -822 291747 299134 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 4913 298990 5223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 13913 298990 14223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 22913 298990 23223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 31913 298990 32223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 40913 298990 41223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 49913 298990 50223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 58913 298990 59223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 67913 298990 68223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 76913 298990 77223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 85913 298990 86223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 94913 298990 95223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 103913 298990 104223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 112913 298990 113223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 121913 298990 122223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 130913 298990 131223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 139913 298990 140223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 148913 298990 149223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 157913 298990 158223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 166913 298990 167223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 175913 298990 176223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 184913 298990 185223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 193913 298990 194223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 202913 298990 203223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 211913 298990 212223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 220913 298990 221223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 229913 298990 230223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 238913 298990 239223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 247913 298990 248223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 256913 298990 257223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 265913 298990 266223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 274913 298990 275223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 283913 298990 284223 6 vss
port 533 nsew ground bidirectional
rlabel metal5 s -958 292913 298990 293223 6 vss
port 533 nsew ground bidirectional
rlabel metal2 s 10892 -480 11004 240 8 wb_clk_i
port 534 nsew signal input
rlabel metal2 s 11452 -480 11564 240 8 wb_rst_i
port 535 nsew signal input
rlabel metal2 s 12012 -480 12124 240 8 wbs_ack_o
port 536 nsew signal output
rlabel metal2 s 14252 -480 14364 240 8 wbs_adr_i[0]
port 537 nsew signal input
rlabel metal2 s 33292 -480 33404 240 8 wbs_adr_i[10]
port 538 nsew signal input
rlabel metal2 s 34972 -480 35084 240 8 wbs_adr_i[11]
port 539 nsew signal input
rlabel metal2 s 36652 -480 36764 240 8 wbs_adr_i[12]
port 540 nsew signal input
rlabel metal2 s 38332 -480 38444 240 8 wbs_adr_i[13]
port 541 nsew signal input
rlabel metal2 s 40012 -480 40124 240 8 wbs_adr_i[14]
port 542 nsew signal input
rlabel metal2 s 41692 -480 41804 240 8 wbs_adr_i[15]
port 543 nsew signal input
rlabel metal2 s 43372 -480 43484 240 8 wbs_adr_i[16]
port 544 nsew signal input
rlabel metal2 s 45052 -480 45164 240 8 wbs_adr_i[17]
port 545 nsew signal input
rlabel metal2 s 46732 -480 46844 240 8 wbs_adr_i[18]
port 546 nsew signal input
rlabel metal2 s 48412 -480 48524 240 8 wbs_adr_i[19]
port 547 nsew signal input
rlabel metal2 s 16492 -480 16604 240 8 wbs_adr_i[1]
port 548 nsew signal input
rlabel metal2 s 50092 -480 50204 240 8 wbs_adr_i[20]
port 549 nsew signal input
rlabel metal2 s 51772 -480 51884 240 8 wbs_adr_i[21]
port 550 nsew signal input
rlabel metal2 s 53452 -480 53564 240 8 wbs_adr_i[22]
port 551 nsew signal input
rlabel metal2 s 55132 -480 55244 240 8 wbs_adr_i[23]
port 552 nsew signal input
rlabel metal2 s 56812 -480 56924 240 8 wbs_adr_i[24]
port 553 nsew signal input
rlabel metal2 s 58492 -480 58604 240 8 wbs_adr_i[25]
port 554 nsew signal input
rlabel metal2 s 60172 -480 60284 240 8 wbs_adr_i[26]
port 555 nsew signal input
rlabel metal2 s 61852 -480 61964 240 8 wbs_adr_i[27]
port 556 nsew signal input
rlabel metal2 s 63532 -480 63644 240 8 wbs_adr_i[28]
port 557 nsew signal input
rlabel metal2 s 65212 -480 65324 240 8 wbs_adr_i[29]
port 558 nsew signal input
rlabel metal2 s 18732 -480 18844 240 8 wbs_adr_i[2]
port 559 nsew signal input
rlabel metal2 s 66892 -480 67004 240 8 wbs_adr_i[30]
port 560 nsew signal input
rlabel metal2 s 68572 -480 68684 240 8 wbs_adr_i[31]
port 561 nsew signal input
rlabel metal2 s 20972 -480 21084 240 8 wbs_adr_i[3]
port 562 nsew signal input
rlabel metal2 s 23212 -480 23324 240 8 wbs_adr_i[4]
port 563 nsew signal input
rlabel metal2 s 24892 -480 25004 240 8 wbs_adr_i[5]
port 564 nsew signal input
rlabel metal2 s 26572 -480 26684 240 8 wbs_adr_i[6]
port 565 nsew signal input
rlabel metal2 s 28252 -480 28364 240 8 wbs_adr_i[7]
port 566 nsew signal input
rlabel metal2 s 29932 -480 30044 240 8 wbs_adr_i[8]
port 567 nsew signal input
rlabel metal2 s 31612 -480 31724 240 8 wbs_adr_i[9]
port 568 nsew signal input
rlabel metal2 s 12572 -480 12684 240 8 wbs_cyc_i
port 569 nsew signal input
rlabel metal2 s 14812 -480 14924 240 8 wbs_dat_i[0]
port 570 nsew signal input
rlabel metal2 s 33852 -480 33964 240 8 wbs_dat_i[10]
port 571 nsew signal input
rlabel metal2 s 35532 -480 35644 240 8 wbs_dat_i[11]
port 572 nsew signal input
rlabel metal2 s 37212 -480 37324 240 8 wbs_dat_i[12]
port 573 nsew signal input
rlabel metal2 s 38892 -480 39004 240 8 wbs_dat_i[13]
port 574 nsew signal input
rlabel metal2 s 40572 -480 40684 240 8 wbs_dat_i[14]
port 575 nsew signal input
rlabel metal2 s 42252 -480 42364 240 8 wbs_dat_i[15]
port 576 nsew signal input
rlabel metal2 s 43932 -480 44044 240 8 wbs_dat_i[16]
port 577 nsew signal input
rlabel metal2 s 45612 -480 45724 240 8 wbs_dat_i[17]
port 578 nsew signal input
rlabel metal2 s 47292 -480 47404 240 8 wbs_dat_i[18]
port 579 nsew signal input
rlabel metal2 s 48972 -480 49084 240 8 wbs_dat_i[19]
port 580 nsew signal input
rlabel metal2 s 17052 -480 17164 240 8 wbs_dat_i[1]
port 581 nsew signal input
rlabel metal2 s 50652 -480 50764 240 8 wbs_dat_i[20]
port 582 nsew signal input
rlabel metal2 s 52332 -480 52444 240 8 wbs_dat_i[21]
port 583 nsew signal input
rlabel metal2 s 54012 -480 54124 240 8 wbs_dat_i[22]
port 584 nsew signal input
rlabel metal2 s 55692 -480 55804 240 8 wbs_dat_i[23]
port 585 nsew signal input
rlabel metal2 s 57372 -480 57484 240 8 wbs_dat_i[24]
port 586 nsew signal input
rlabel metal2 s 59052 -480 59164 240 8 wbs_dat_i[25]
port 587 nsew signal input
rlabel metal2 s 60732 -480 60844 240 8 wbs_dat_i[26]
port 588 nsew signal input
rlabel metal2 s 62412 -480 62524 240 8 wbs_dat_i[27]
port 589 nsew signal input
rlabel metal2 s 64092 -480 64204 240 8 wbs_dat_i[28]
port 590 nsew signal input
rlabel metal2 s 65772 -480 65884 240 8 wbs_dat_i[29]
port 591 nsew signal input
rlabel metal2 s 19292 -480 19404 240 8 wbs_dat_i[2]
port 592 nsew signal input
rlabel metal2 s 67452 -480 67564 240 8 wbs_dat_i[30]
port 593 nsew signal input
rlabel metal2 s 69132 -480 69244 240 8 wbs_dat_i[31]
port 594 nsew signal input
rlabel metal2 s 21532 -480 21644 240 8 wbs_dat_i[3]
port 595 nsew signal input
rlabel metal2 s 23772 -480 23884 240 8 wbs_dat_i[4]
port 596 nsew signal input
rlabel metal2 s 25452 -480 25564 240 8 wbs_dat_i[5]
port 597 nsew signal input
rlabel metal2 s 27132 -480 27244 240 8 wbs_dat_i[6]
port 598 nsew signal input
rlabel metal2 s 28812 -480 28924 240 8 wbs_dat_i[7]
port 599 nsew signal input
rlabel metal2 s 30492 -480 30604 240 8 wbs_dat_i[8]
port 600 nsew signal input
rlabel metal2 s 32172 -480 32284 240 8 wbs_dat_i[9]
port 601 nsew signal input
rlabel metal2 s 15372 -480 15484 240 8 wbs_dat_o[0]
port 602 nsew signal output
rlabel metal2 s 34412 -480 34524 240 8 wbs_dat_o[10]
port 603 nsew signal output
rlabel metal2 s 36092 -480 36204 240 8 wbs_dat_o[11]
port 604 nsew signal output
rlabel metal2 s 37772 -480 37884 240 8 wbs_dat_o[12]
port 605 nsew signal output
rlabel metal2 s 39452 -480 39564 240 8 wbs_dat_o[13]
port 606 nsew signal output
rlabel metal2 s 41132 -480 41244 240 8 wbs_dat_o[14]
port 607 nsew signal output
rlabel metal2 s 42812 -480 42924 240 8 wbs_dat_o[15]
port 608 nsew signal output
rlabel metal2 s 44492 -480 44604 240 8 wbs_dat_o[16]
port 609 nsew signal output
rlabel metal2 s 46172 -480 46284 240 8 wbs_dat_o[17]
port 610 nsew signal output
rlabel metal2 s 47852 -480 47964 240 8 wbs_dat_o[18]
port 611 nsew signal output
rlabel metal2 s 49532 -480 49644 240 8 wbs_dat_o[19]
port 612 nsew signal output
rlabel metal2 s 17612 -480 17724 240 8 wbs_dat_o[1]
port 613 nsew signal output
rlabel metal2 s 51212 -480 51324 240 8 wbs_dat_o[20]
port 614 nsew signal output
rlabel metal2 s 52892 -480 53004 240 8 wbs_dat_o[21]
port 615 nsew signal output
rlabel metal2 s 54572 -480 54684 240 8 wbs_dat_o[22]
port 616 nsew signal output
rlabel metal2 s 56252 -480 56364 240 8 wbs_dat_o[23]
port 617 nsew signal output
rlabel metal2 s 57932 -480 58044 240 8 wbs_dat_o[24]
port 618 nsew signal output
rlabel metal2 s 59612 -480 59724 240 8 wbs_dat_o[25]
port 619 nsew signal output
rlabel metal2 s 61292 -480 61404 240 8 wbs_dat_o[26]
port 620 nsew signal output
rlabel metal2 s 62972 -480 63084 240 8 wbs_dat_o[27]
port 621 nsew signal output
rlabel metal2 s 64652 -480 64764 240 8 wbs_dat_o[28]
port 622 nsew signal output
rlabel metal2 s 66332 -480 66444 240 8 wbs_dat_o[29]
port 623 nsew signal output
rlabel metal2 s 19852 -480 19964 240 8 wbs_dat_o[2]
port 624 nsew signal output
rlabel metal2 s 68012 -480 68124 240 8 wbs_dat_o[30]
port 625 nsew signal output
rlabel metal2 s 69692 -480 69804 240 8 wbs_dat_o[31]
port 626 nsew signal output
rlabel metal2 s 22092 -480 22204 240 8 wbs_dat_o[3]
port 627 nsew signal output
rlabel metal2 s 24332 -480 24444 240 8 wbs_dat_o[4]
port 628 nsew signal output
rlabel metal2 s 26012 -480 26124 240 8 wbs_dat_o[5]
port 629 nsew signal output
rlabel metal2 s 27692 -480 27804 240 8 wbs_dat_o[6]
port 630 nsew signal output
rlabel metal2 s 29372 -480 29484 240 8 wbs_dat_o[7]
port 631 nsew signal output
rlabel metal2 s 31052 -480 31164 240 8 wbs_dat_o[8]
port 632 nsew signal output
rlabel metal2 s 32732 -480 32844 240 8 wbs_dat_o[9]
port 633 nsew signal output
rlabel metal2 s 15932 -480 16044 240 8 wbs_sel_i[0]
port 634 nsew signal input
rlabel metal2 s 18172 -480 18284 240 8 wbs_sel_i[1]
port 635 nsew signal input
rlabel metal2 s 20412 -480 20524 240 8 wbs_sel_i[2]
port 636 nsew signal input
rlabel metal2 s 22652 -480 22764 240 8 wbs_sel_i[3]
port 637 nsew signal input
rlabel metal2 s 13132 -480 13244 240 8 wbs_stb_i
port 638 nsew signal input
rlabel metal2 s 13692 -480 13804 240 8 wbs_we_i
port 639 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 298020 298020
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 5706100
string GDS_FILE /opt/caravel_180/openlane/user_project_wrapper/runs/22_12_03_04_07/results/signoff/user_project_wrapper.magic.gds
string GDS_START 2526948
<< end >>

