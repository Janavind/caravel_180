VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO macro_golden
  CLASS BLOCK ;
  FOREIGN macro_golden ;
  ORIGIN 0.000 0.000 ;
  SIZE 600.000 BY 600.000 ;
  PIN io_active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 12.320 596.000 12.880 600.000 ;
    END
  END io_active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 17.360 596.000 17.920 600.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 168.560 596.000 169.120 600.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 183.680 596.000 184.240 600.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 198.800 596.000 199.360 600.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 213.920 596.000 214.480 600.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 229.040 596.000 229.600 600.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 244.160 596.000 244.720 600.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 259.280 596.000 259.840 600.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 274.400 596.000 274.960 600.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 289.520 596.000 290.080 600.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 304.640 596.000 305.200 600.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 32.480 596.000 33.040 600.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 319.760 596.000 320.320 600.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 334.880 596.000 335.440 600.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 350.000 596.000 350.560 600.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 365.120 596.000 365.680 600.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 380.240 596.000 380.800 600.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 395.360 596.000 395.920 600.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 410.480 596.000 411.040 600.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 425.600 596.000 426.160 600.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 440.720 596.000 441.280 600.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 455.840 596.000 456.400 600.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 47.600 596.000 48.160 600.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 470.960 596.000 471.520 600.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 486.080 596.000 486.640 600.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 501.200 596.000 501.760 600.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 516.320 596.000 516.880 600.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 531.440 596.000 532.000 600.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 546.560 596.000 547.120 600.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 561.680 596.000 562.240 600.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 576.800 596.000 577.360 600.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 62.720 596.000 63.280 600.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 77.840 596.000 78.400 600.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 92.960 596.000 93.520 600.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 108.080 596.000 108.640 600.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 123.200 596.000 123.760 600.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 138.320 596.000 138.880 600.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 153.440 596.000 154.000 600.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 22.400 596.000 22.960 600.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 173.600 596.000 174.160 600.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 188.720 596.000 189.280 600.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 203.840 596.000 204.400 600.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 218.960 596.000 219.520 600.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 234.080 596.000 234.640 600.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 249.200 596.000 249.760 600.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 264.320 596.000 264.880 600.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 279.440 596.000 280.000 600.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 294.560 596.000 295.120 600.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 309.680 596.000 310.240 600.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 37.520 596.000 38.080 600.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 324.800 596.000 325.360 600.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 339.920 596.000 340.480 600.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 355.040 596.000 355.600 600.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 370.160 596.000 370.720 600.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 385.280 596.000 385.840 600.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 400.400 596.000 400.960 600.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 415.520 596.000 416.080 600.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 430.640 596.000 431.200 600.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 445.760 596.000 446.320 600.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 460.880 596.000 461.440 600.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 52.640 596.000 53.200 600.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 476.000 596.000 476.560 600.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 491.120 596.000 491.680 600.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 506.240 596.000 506.800 600.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 521.360 596.000 521.920 600.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 536.480 596.000 537.040 600.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 551.600 596.000 552.160 600.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 566.720 596.000 567.280 600.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 581.840 596.000 582.400 600.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 67.760 596.000 68.320 600.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 82.880 596.000 83.440 600.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 98.000 596.000 98.560 600.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 113.120 596.000 113.680 600.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 128.240 596.000 128.800 600.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 143.360 596.000 143.920 600.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 158.480 596.000 159.040 600.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 27.440 596.000 28.000 600.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 178.640 596.000 179.200 600.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 193.760 596.000 194.320 600.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 208.880 596.000 209.440 600.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 224.000 596.000 224.560 600.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 239.120 596.000 239.680 600.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 254.240 596.000 254.800 600.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 269.360 596.000 269.920 600.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 284.480 596.000 285.040 600.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 299.600 596.000 300.160 600.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 314.720 596.000 315.280 600.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 42.560 596.000 43.120 600.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 329.840 596.000 330.400 600.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 344.960 596.000 345.520 600.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 360.080 596.000 360.640 600.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 375.200 596.000 375.760 600.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 390.320 596.000 390.880 600.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 405.440 596.000 406.000 600.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 420.560 596.000 421.120 600.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 435.680 596.000 436.240 600.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 450.800 596.000 451.360 600.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 465.920 596.000 466.480 600.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 57.680 596.000 58.240 600.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 481.040 596.000 481.600 600.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 496.160 596.000 496.720 600.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 511.280 596.000 511.840 600.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 526.400 596.000 526.960 600.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 541.520 596.000 542.080 600.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 556.640 596.000 557.200 600.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 571.760 596.000 572.320 600.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 586.880 596.000 587.440 600.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 72.800 596.000 73.360 600.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 87.920 596.000 88.480 600.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 103.040 596.000 103.600 600.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 118.160 596.000 118.720 600.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 133.280 596.000 133.840 600.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 148.400 596.000 148.960 600.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 163.520 596.000 164.080 600.000 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 227.920 0.000 228.480 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 278.320 0.000 278.880 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 283.360 0.000 283.920 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 288.400 0.000 288.960 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 293.440 0.000 294.000 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 298.480 0.000 299.040 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 303.520 0.000 304.080 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 308.560 0.000 309.120 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 313.600 0.000 314.160 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 318.640 0.000 319.200 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 323.680 0.000 324.240 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 232.960 0.000 233.520 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 328.720 0.000 329.280 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 333.760 0.000 334.320 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 338.800 0.000 339.360 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 343.840 0.000 344.400 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 348.880 0.000 349.440 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 353.920 0.000 354.480 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 358.960 0.000 359.520 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 364.000 0.000 364.560 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 369.040 0.000 369.600 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 374.080 0.000 374.640 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 238.000 0.000 238.560 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 379.120 0.000 379.680 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 384.160 0.000 384.720 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 389.200 0.000 389.760 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 394.240 0.000 394.800 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 399.280 0.000 399.840 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 404.320 0.000 404.880 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 409.360 0.000 409.920 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 414.400 0.000 414.960 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 419.440 0.000 420.000 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 424.480 0.000 425.040 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 243.040 0.000 243.600 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 429.520 0.000 430.080 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 434.560 0.000 435.120 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 439.600 0.000 440.160 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 444.640 0.000 445.200 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 449.680 0.000 450.240 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 454.720 0.000 455.280 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 459.760 0.000 460.320 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 464.800 0.000 465.360 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 469.840 0.000 470.400 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 474.880 0.000 475.440 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 248.080 0.000 248.640 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 479.920 0.000 480.480 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 484.960 0.000 485.520 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 490.000 0.000 490.560 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 495.040 0.000 495.600 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 500.080 0.000 500.640 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 505.120 0.000 505.680 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 510.160 0.000 510.720 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 515.200 0.000 515.760 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 520.240 0.000 520.800 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 525.280 0.000 525.840 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 253.120 0.000 253.680 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 530.320 0.000 530.880 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 535.360 0.000 535.920 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 540.400 0.000 540.960 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 545.440 0.000 546.000 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 258.160 0.000 258.720 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 263.200 0.000 263.760 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 268.240 0.000 268.800 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 273.280 0.000 273.840 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 229.600 0.000 230.160 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 280.000 0.000 280.560 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 285.040 0.000 285.600 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 290.080 0.000 290.640 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 295.120 0.000 295.680 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 300.160 0.000 300.720 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 305.200 0.000 305.760 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 310.240 0.000 310.800 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 315.280 0.000 315.840 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 320.320 0.000 320.880 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 325.360 0.000 325.920 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 234.640 0.000 235.200 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 330.400 0.000 330.960 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 335.440 0.000 336.000 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 340.480 0.000 341.040 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 345.520 0.000 346.080 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 350.560 0.000 351.120 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 355.600 0.000 356.160 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 360.640 0.000 361.200 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 365.680 0.000 366.240 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 370.720 0.000 371.280 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 375.760 0.000 376.320 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 239.680 0.000 240.240 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 380.800 0.000 381.360 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 385.840 0.000 386.400 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 390.880 0.000 391.440 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 395.920 0.000 396.480 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 400.960 0.000 401.520 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 406.000 0.000 406.560 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 411.040 0.000 411.600 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 416.080 0.000 416.640 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 421.120 0.000 421.680 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 426.160 0.000 426.720 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 244.720 0.000 245.280 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 431.200 0.000 431.760 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 436.240 0.000 436.800 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 441.280 0.000 441.840 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 446.320 0.000 446.880 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 451.360 0.000 451.920 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 456.400 0.000 456.960 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 461.440 0.000 462.000 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 466.480 0.000 467.040 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 471.520 0.000 472.080 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 476.560 0.000 477.120 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 249.760 0.000 250.320 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 481.600 0.000 482.160 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 486.640 0.000 487.200 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 491.680 0.000 492.240 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 496.720 0.000 497.280 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 501.760 0.000 502.320 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 506.800 0.000 507.360 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 511.840 0.000 512.400 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 516.880 0.000 517.440 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 521.920 0.000 522.480 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 526.960 0.000 527.520 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 254.800 0.000 255.360 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 532.000 0.000 532.560 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 537.040 0.000 537.600 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 542.080 0.000 542.640 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 547.120 0.000 547.680 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 259.840 0.000 260.400 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 264.880 0.000 265.440 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 269.920 0.000 270.480 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 274.960 0.000 275.520 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 231.280 0.000 231.840 4.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 281.680 0.000 282.240 4.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 286.720 0.000 287.280 4.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 291.760 0.000 292.320 4.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 296.800 0.000 297.360 4.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 301.840 0.000 302.400 4.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 306.880 0.000 307.440 4.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 311.920 0.000 312.480 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 316.960 0.000 317.520 4.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 322.000 0.000 322.560 4.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 327.040 0.000 327.600 4.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 236.320 0.000 236.880 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 332.080 0.000 332.640 4.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 337.120 0.000 337.680 4.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 342.160 0.000 342.720 4.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 347.200 0.000 347.760 4.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 352.240 0.000 352.800 4.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 357.280 0.000 357.840 4.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 362.320 0.000 362.880 4.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 367.360 0.000 367.920 4.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 372.400 0.000 372.960 4.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 377.440 0.000 378.000 4.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 241.360 0.000 241.920 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 382.480 0.000 383.040 4.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 387.520 0.000 388.080 4.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 392.560 0.000 393.120 4.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 397.600 0.000 398.160 4.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 402.640 0.000 403.200 4.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 407.680 0.000 408.240 4.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 412.720 0.000 413.280 4.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 417.760 0.000 418.320 4.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 422.800 0.000 423.360 4.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 427.840 0.000 428.400 4.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 246.400 0.000 246.960 4.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 432.880 0.000 433.440 4.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 437.920 0.000 438.480 4.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 442.960 0.000 443.520 4.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 448.000 0.000 448.560 4.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 453.040 0.000 453.600 4.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 458.080 0.000 458.640 4.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 463.120 0.000 463.680 4.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 468.160 0.000 468.720 4.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 473.200 0.000 473.760 4.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 478.240 0.000 478.800 4.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 251.440 0.000 252.000 4.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 483.280 0.000 483.840 4.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 488.320 0.000 488.880 4.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 493.360 0.000 493.920 4.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 498.400 0.000 498.960 4.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 503.440 0.000 504.000 4.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 508.480 0.000 509.040 4.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 513.520 0.000 514.080 4.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 518.560 0.000 519.120 4.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 523.600 0.000 524.160 4.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 528.640 0.000 529.200 4.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 256.480 0.000 257.040 4.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 533.680 0.000 534.240 4.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 538.720 0.000 539.280 4.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 543.760 0.000 544.320 4.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 548.800 0.000 549.360 4.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 261.520 0.000 262.080 4.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 266.560 0.000 267.120 4.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 271.600 0.000 272.160 4.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 276.640 0.000 277.200 4.000 ;
    END
  END la_oenb[9]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 584.380 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 584.380 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 49.840 0.000 50.400 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 51.520 0.000 52.080 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 53.200 0.000 53.760 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 59.920 0.000 60.480 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 117.040 0.000 117.600 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 122.080 0.000 122.640 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 127.120 0.000 127.680 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 132.160 0.000 132.720 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 137.200 0.000 137.760 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 142.240 0.000 142.800 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 147.280 0.000 147.840 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 152.320 0.000 152.880 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 157.360 0.000 157.920 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 162.400 0.000 162.960 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 66.640 0.000 67.200 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 167.440 0.000 168.000 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 172.480 0.000 173.040 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 177.520 0.000 178.080 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 182.560 0.000 183.120 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 187.600 0.000 188.160 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 192.640 0.000 193.200 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 197.680 0.000 198.240 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 202.720 0.000 203.280 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 207.760 0.000 208.320 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 212.800 0.000 213.360 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 73.360 0.000 73.920 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 217.840 0.000 218.400 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 222.880 0.000 223.440 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 80.080 0.000 80.640 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 86.800 0.000 87.360 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 91.840 0.000 92.400 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 96.880 0.000 97.440 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 101.920 0.000 102.480 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 106.960 0.000 107.520 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 112.000 0.000 112.560 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 54.880 0.000 55.440 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 61.600 0.000 62.160 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 118.720 0.000 119.280 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 123.760 0.000 124.320 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 128.800 0.000 129.360 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 133.840 0.000 134.400 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 138.880 0.000 139.440 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 143.920 0.000 144.480 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 148.960 0.000 149.520 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 154.000 0.000 154.560 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 159.040 0.000 159.600 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 164.080 0.000 164.640 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 68.320 0.000 68.880 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 169.120 0.000 169.680 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 174.160 0.000 174.720 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 179.200 0.000 179.760 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 184.240 0.000 184.800 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 189.280 0.000 189.840 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 194.320 0.000 194.880 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 199.360 0.000 199.920 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 204.400 0.000 204.960 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 209.440 0.000 210.000 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 214.480 0.000 215.040 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 75.040 0.000 75.600 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 219.520 0.000 220.080 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 224.560 0.000 225.120 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 81.760 0.000 82.320 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 88.480 0.000 89.040 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 93.520 0.000 94.080 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 98.560 0.000 99.120 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 103.600 0.000 104.160 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 108.640 0.000 109.200 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 113.680 0.000 114.240 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 63.280 0.000 63.840 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 120.400 0.000 120.960 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 125.440 0.000 126.000 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 130.480 0.000 131.040 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 135.520 0.000 136.080 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 140.560 0.000 141.120 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 145.600 0.000 146.160 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 150.640 0.000 151.200 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 155.680 0.000 156.240 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 160.720 0.000 161.280 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 165.760 0.000 166.320 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 70.000 0.000 70.560 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 170.800 0.000 171.360 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 175.840 0.000 176.400 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 180.880 0.000 181.440 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 185.920 0.000 186.480 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 190.960 0.000 191.520 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 196.000 0.000 196.560 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 201.040 0.000 201.600 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 206.080 0.000 206.640 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 211.120 0.000 211.680 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 216.160 0.000 216.720 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 76.720 0.000 77.280 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 221.200 0.000 221.760 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 226.240 0.000 226.800 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 83.440 0.000 84.000 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 90.160 0.000 90.720 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 95.200 0.000 95.760 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 100.240 0.000 100.800 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 105.280 0.000 105.840 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 110.320 0.000 110.880 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 115.360 0.000 115.920 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 64.960 0.000 65.520 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 71.680 0.000 72.240 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 78.400 0.000 78.960 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 85.120 0.000 85.680 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 56.560 0.000 57.120 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 58.240 0.000 58.800 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 8.550 593.040 586.730 ;
      LAYER Metal2 ;
        RECT 11.340 595.700 12.020 596.820 ;
        RECT 13.180 595.700 17.060 596.820 ;
        RECT 18.220 595.700 22.100 596.820 ;
        RECT 23.260 595.700 27.140 596.820 ;
        RECT 28.300 595.700 32.180 596.820 ;
        RECT 33.340 595.700 37.220 596.820 ;
        RECT 38.380 595.700 42.260 596.820 ;
        RECT 43.420 595.700 47.300 596.820 ;
        RECT 48.460 595.700 52.340 596.820 ;
        RECT 53.500 595.700 57.380 596.820 ;
        RECT 58.540 595.700 62.420 596.820 ;
        RECT 63.580 595.700 67.460 596.820 ;
        RECT 68.620 595.700 72.500 596.820 ;
        RECT 73.660 595.700 77.540 596.820 ;
        RECT 78.700 595.700 82.580 596.820 ;
        RECT 83.740 595.700 87.620 596.820 ;
        RECT 88.780 595.700 92.660 596.820 ;
        RECT 93.820 595.700 97.700 596.820 ;
        RECT 98.860 595.700 102.740 596.820 ;
        RECT 103.900 595.700 107.780 596.820 ;
        RECT 108.940 595.700 112.820 596.820 ;
        RECT 113.980 595.700 117.860 596.820 ;
        RECT 119.020 595.700 122.900 596.820 ;
        RECT 124.060 595.700 127.940 596.820 ;
        RECT 129.100 595.700 132.980 596.820 ;
        RECT 134.140 595.700 138.020 596.820 ;
        RECT 139.180 595.700 143.060 596.820 ;
        RECT 144.220 595.700 148.100 596.820 ;
        RECT 149.260 595.700 153.140 596.820 ;
        RECT 154.300 595.700 158.180 596.820 ;
        RECT 159.340 595.700 163.220 596.820 ;
        RECT 164.380 595.700 168.260 596.820 ;
        RECT 169.420 595.700 173.300 596.820 ;
        RECT 174.460 595.700 178.340 596.820 ;
        RECT 179.500 595.700 183.380 596.820 ;
        RECT 184.540 595.700 188.420 596.820 ;
        RECT 189.580 595.700 193.460 596.820 ;
        RECT 194.620 595.700 198.500 596.820 ;
        RECT 199.660 595.700 203.540 596.820 ;
        RECT 204.700 595.700 208.580 596.820 ;
        RECT 209.740 595.700 213.620 596.820 ;
        RECT 214.780 595.700 218.660 596.820 ;
        RECT 219.820 595.700 223.700 596.820 ;
        RECT 224.860 595.700 228.740 596.820 ;
        RECT 229.900 595.700 233.780 596.820 ;
        RECT 234.940 595.700 238.820 596.820 ;
        RECT 239.980 595.700 243.860 596.820 ;
        RECT 245.020 595.700 248.900 596.820 ;
        RECT 250.060 595.700 253.940 596.820 ;
        RECT 255.100 595.700 258.980 596.820 ;
        RECT 260.140 595.700 264.020 596.820 ;
        RECT 265.180 595.700 269.060 596.820 ;
        RECT 270.220 595.700 274.100 596.820 ;
        RECT 275.260 595.700 279.140 596.820 ;
        RECT 280.300 595.700 284.180 596.820 ;
        RECT 285.340 595.700 289.220 596.820 ;
        RECT 290.380 595.700 294.260 596.820 ;
        RECT 295.420 595.700 299.300 596.820 ;
        RECT 300.460 595.700 304.340 596.820 ;
        RECT 305.500 595.700 309.380 596.820 ;
        RECT 310.540 595.700 314.420 596.820 ;
        RECT 315.580 595.700 319.460 596.820 ;
        RECT 320.620 595.700 324.500 596.820 ;
        RECT 325.660 595.700 329.540 596.820 ;
        RECT 330.700 595.700 334.580 596.820 ;
        RECT 335.740 595.700 339.620 596.820 ;
        RECT 340.780 595.700 344.660 596.820 ;
        RECT 345.820 595.700 349.700 596.820 ;
        RECT 350.860 595.700 354.740 596.820 ;
        RECT 355.900 595.700 359.780 596.820 ;
        RECT 360.940 595.700 364.820 596.820 ;
        RECT 365.980 595.700 369.860 596.820 ;
        RECT 371.020 595.700 374.900 596.820 ;
        RECT 376.060 595.700 379.940 596.820 ;
        RECT 381.100 595.700 384.980 596.820 ;
        RECT 386.140 595.700 390.020 596.820 ;
        RECT 391.180 595.700 395.060 596.820 ;
        RECT 396.220 595.700 400.100 596.820 ;
        RECT 401.260 595.700 405.140 596.820 ;
        RECT 406.300 595.700 410.180 596.820 ;
        RECT 411.340 595.700 415.220 596.820 ;
        RECT 416.380 595.700 420.260 596.820 ;
        RECT 421.420 595.700 425.300 596.820 ;
        RECT 426.460 595.700 430.340 596.820 ;
        RECT 431.500 595.700 435.380 596.820 ;
        RECT 436.540 595.700 440.420 596.820 ;
        RECT 441.580 595.700 445.460 596.820 ;
        RECT 446.620 595.700 450.500 596.820 ;
        RECT 451.660 595.700 455.540 596.820 ;
        RECT 456.700 595.700 460.580 596.820 ;
        RECT 461.740 595.700 465.620 596.820 ;
        RECT 466.780 595.700 470.660 596.820 ;
        RECT 471.820 595.700 475.700 596.820 ;
        RECT 476.860 595.700 480.740 596.820 ;
        RECT 481.900 595.700 485.780 596.820 ;
        RECT 486.940 595.700 490.820 596.820 ;
        RECT 491.980 595.700 495.860 596.820 ;
        RECT 497.020 595.700 500.900 596.820 ;
        RECT 502.060 595.700 505.940 596.820 ;
        RECT 507.100 595.700 510.980 596.820 ;
        RECT 512.140 595.700 516.020 596.820 ;
        RECT 517.180 595.700 521.060 596.820 ;
        RECT 522.220 595.700 526.100 596.820 ;
        RECT 527.260 595.700 531.140 596.820 ;
        RECT 532.300 595.700 536.180 596.820 ;
        RECT 537.340 595.700 541.220 596.820 ;
        RECT 542.380 595.700 546.260 596.820 ;
        RECT 547.420 595.700 551.300 596.820 ;
        RECT 552.460 595.700 556.340 596.820 ;
        RECT 557.500 595.700 561.380 596.820 ;
        RECT 562.540 595.700 566.420 596.820 ;
        RECT 567.580 595.700 571.460 596.820 ;
        RECT 572.620 595.700 576.500 596.820 ;
        RECT 577.660 595.700 581.540 596.820 ;
        RECT 582.700 595.700 586.580 596.820 ;
        RECT 587.740 595.700 588.420 596.820 ;
        RECT 11.340 4.300 588.420 595.700 ;
        RECT 11.340 4.000 49.540 4.300 ;
        RECT 50.700 4.000 51.220 4.300 ;
        RECT 52.380 4.000 52.900 4.300 ;
        RECT 54.060 4.000 54.580 4.300 ;
        RECT 55.740 4.000 56.260 4.300 ;
        RECT 57.420 4.000 57.940 4.300 ;
        RECT 59.100 4.000 59.620 4.300 ;
        RECT 60.780 4.000 61.300 4.300 ;
        RECT 62.460 4.000 62.980 4.300 ;
        RECT 64.140 4.000 64.660 4.300 ;
        RECT 65.820 4.000 66.340 4.300 ;
        RECT 67.500 4.000 68.020 4.300 ;
        RECT 69.180 4.000 69.700 4.300 ;
        RECT 70.860 4.000 71.380 4.300 ;
        RECT 72.540 4.000 73.060 4.300 ;
        RECT 74.220 4.000 74.740 4.300 ;
        RECT 75.900 4.000 76.420 4.300 ;
        RECT 77.580 4.000 78.100 4.300 ;
        RECT 79.260 4.000 79.780 4.300 ;
        RECT 80.940 4.000 81.460 4.300 ;
        RECT 82.620 4.000 83.140 4.300 ;
        RECT 84.300 4.000 84.820 4.300 ;
        RECT 85.980 4.000 86.500 4.300 ;
        RECT 87.660 4.000 88.180 4.300 ;
        RECT 89.340 4.000 89.860 4.300 ;
        RECT 91.020 4.000 91.540 4.300 ;
        RECT 92.700 4.000 93.220 4.300 ;
        RECT 94.380 4.000 94.900 4.300 ;
        RECT 96.060 4.000 96.580 4.300 ;
        RECT 97.740 4.000 98.260 4.300 ;
        RECT 99.420 4.000 99.940 4.300 ;
        RECT 101.100 4.000 101.620 4.300 ;
        RECT 102.780 4.000 103.300 4.300 ;
        RECT 104.460 4.000 104.980 4.300 ;
        RECT 106.140 4.000 106.660 4.300 ;
        RECT 107.820 4.000 108.340 4.300 ;
        RECT 109.500 4.000 110.020 4.300 ;
        RECT 111.180 4.000 111.700 4.300 ;
        RECT 112.860 4.000 113.380 4.300 ;
        RECT 114.540 4.000 115.060 4.300 ;
        RECT 116.220 4.000 116.740 4.300 ;
        RECT 117.900 4.000 118.420 4.300 ;
        RECT 119.580 4.000 120.100 4.300 ;
        RECT 121.260 4.000 121.780 4.300 ;
        RECT 122.940 4.000 123.460 4.300 ;
        RECT 124.620 4.000 125.140 4.300 ;
        RECT 126.300 4.000 126.820 4.300 ;
        RECT 127.980 4.000 128.500 4.300 ;
        RECT 129.660 4.000 130.180 4.300 ;
        RECT 131.340 4.000 131.860 4.300 ;
        RECT 133.020 4.000 133.540 4.300 ;
        RECT 134.700 4.000 135.220 4.300 ;
        RECT 136.380 4.000 136.900 4.300 ;
        RECT 138.060 4.000 138.580 4.300 ;
        RECT 139.740 4.000 140.260 4.300 ;
        RECT 141.420 4.000 141.940 4.300 ;
        RECT 143.100 4.000 143.620 4.300 ;
        RECT 144.780 4.000 145.300 4.300 ;
        RECT 146.460 4.000 146.980 4.300 ;
        RECT 148.140 4.000 148.660 4.300 ;
        RECT 149.820 4.000 150.340 4.300 ;
        RECT 151.500 4.000 152.020 4.300 ;
        RECT 153.180 4.000 153.700 4.300 ;
        RECT 154.860 4.000 155.380 4.300 ;
        RECT 156.540 4.000 157.060 4.300 ;
        RECT 158.220 4.000 158.740 4.300 ;
        RECT 159.900 4.000 160.420 4.300 ;
        RECT 161.580 4.000 162.100 4.300 ;
        RECT 163.260 4.000 163.780 4.300 ;
        RECT 164.940 4.000 165.460 4.300 ;
        RECT 166.620 4.000 167.140 4.300 ;
        RECT 168.300 4.000 168.820 4.300 ;
        RECT 169.980 4.000 170.500 4.300 ;
        RECT 171.660 4.000 172.180 4.300 ;
        RECT 173.340 4.000 173.860 4.300 ;
        RECT 175.020 4.000 175.540 4.300 ;
        RECT 176.700 4.000 177.220 4.300 ;
        RECT 178.380 4.000 178.900 4.300 ;
        RECT 180.060 4.000 180.580 4.300 ;
        RECT 181.740 4.000 182.260 4.300 ;
        RECT 183.420 4.000 183.940 4.300 ;
        RECT 185.100 4.000 185.620 4.300 ;
        RECT 186.780 4.000 187.300 4.300 ;
        RECT 188.460 4.000 188.980 4.300 ;
        RECT 190.140 4.000 190.660 4.300 ;
        RECT 191.820 4.000 192.340 4.300 ;
        RECT 193.500 4.000 194.020 4.300 ;
        RECT 195.180 4.000 195.700 4.300 ;
        RECT 196.860 4.000 197.380 4.300 ;
        RECT 198.540 4.000 199.060 4.300 ;
        RECT 200.220 4.000 200.740 4.300 ;
        RECT 201.900 4.000 202.420 4.300 ;
        RECT 203.580 4.000 204.100 4.300 ;
        RECT 205.260 4.000 205.780 4.300 ;
        RECT 206.940 4.000 207.460 4.300 ;
        RECT 208.620 4.000 209.140 4.300 ;
        RECT 210.300 4.000 210.820 4.300 ;
        RECT 211.980 4.000 212.500 4.300 ;
        RECT 213.660 4.000 214.180 4.300 ;
        RECT 215.340 4.000 215.860 4.300 ;
        RECT 217.020 4.000 217.540 4.300 ;
        RECT 218.700 4.000 219.220 4.300 ;
        RECT 220.380 4.000 220.900 4.300 ;
        RECT 222.060 4.000 222.580 4.300 ;
        RECT 223.740 4.000 224.260 4.300 ;
        RECT 225.420 4.000 225.940 4.300 ;
        RECT 227.100 4.000 227.620 4.300 ;
        RECT 228.780 4.000 229.300 4.300 ;
        RECT 230.460 4.000 230.980 4.300 ;
        RECT 232.140 4.000 232.660 4.300 ;
        RECT 233.820 4.000 234.340 4.300 ;
        RECT 235.500 4.000 236.020 4.300 ;
        RECT 237.180 4.000 237.700 4.300 ;
        RECT 238.860 4.000 239.380 4.300 ;
        RECT 240.540 4.000 241.060 4.300 ;
        RECT 242.220 4.000 242.740 4.300 ;
        RECT 243.900 4.000 244.420 4.300 ;
        RECT 245.580 4.000 246.100 4.300 ;
        RECT 247.260 4.000 247.780 4.300 ;
        RECT 248.940 4.000 249.460 4.300 ;
        RECT 250.620 4.000 251.140 4.300 ;
        RECT 252.300 4.000 252.820 4.300 ;
        RECT 253.980 4.000 254.500 4.300 ;
        RECT 255.660 4.000 256.180 4.300 ;
        RECT 257.340 4.000 257.860 4.300 ;
        RECT 259.020 4.000 259.540 4.300 ;
        RECT 260.700 4.000 261.220 4.300 ;
        RECT 262.380 4.000 262.900 4.300 ;
        RECT 264.060 4.000 264.580 4.300 ;
        RECT 265.740 4.000 266.260 4.300 ;
        RECT 267.420 4.000 267.940 4.300 ;
        RECT 269.100 4.000 269.620 4.300 ;
        RECT 270.780 4.000 271.300 4.300 ;
        RECT 272.460 4.000 272.980 4.300 ;
        RECT 274.140 4.000 274.660 4.300 ;
        RECT 275.820 4.000 276.340 4.300 ;
        RECT 277.500 4.000 278.020 4.300 ;
        RECT 279.180 4.000 279.700 4.300 ;
        RECT 280.860 4.000 281.380 4.300 ;
        RECT 282.540 4.000 283.060 4.300 ;
        RECT 284.220 4.000 284.740 4.300 ;
        RECT 285.900 4.000 286.420 4.300 ;
        RECT 287.580 4.000 288.100 4.300 ;
        RECT 289.260 4.000 289.780 4.300 ;
        RECT 290.940 4.000 291.460 4.300 ;
        RECT 292.620 4.000 293.140 4.300 ;
        RECT 294.300 4.000 294.820 4.300 ;
        RECT 295.980 4.000 296.500 4.300 ;
        RECT 297.660 4.000 298.180 4.300 ;
        RECT 299.340 4.000 299.860 4.300 ;
        RECT 301.020 4.000 301.540 4.300 ;
        RECT 302.700 4.000 303.220 4.300 ;
        RECT 304.380 4.000 304.900 4.300 ;
        RECT 306.060 4.000 306.580 4.300 ;
        RECT 307.740 4.000 308.260 4.300 ;
        RECT 309.420 4.000 309.940 4.300 ;
        RECT 311.100 4.000 311.620 4.300 ;
        RECT 312.780 4.000 313.300 4.300 ;
        RECT 314.460 4.000 314.980 4.300 ;
        RECT 316.140 4.000 316.660 4.300 ;
        RECT 317.820 4.000 318.340 4.300 ;
        RECT 319.500 4.000 320.020 4.300 ;
        RECT 321.180 4.000 321.700 4.300 ;
        RECT 322.860 4.000 323.380 4.300 ;
        RECT 324.540 4.000 325.060 4.300 ;
        RECT 326.220 4.000 326.740 4.300 ;
        RECT 327.900 4.000 328.420 4.300 ;
        RECT 329.580 4.000 330.100 4.300 ;
        RECT 331.260 4.000 331.780 4.300 ;
        RECT 332.940 4.000 333.460 4.300 ;
        RECT 334.620 4.000 335.140 4.300 ;
        RECT 336.300 4.000 336.820 4.300 ;
        RECT 337.980 4.000 338.500 4.300 ;
        RECT 339.660 4.000 340.180 4.300 ;
        RECT 341.340 4.000 341.860 4.300 ;
        RECT 343.020 4.000 343.540 4.300 ;
        RECT 344.700 4.000 345.220 4.300 ;
        RECT 346.380 4.000 346.900 4.300 ;
        RECT 348.060 4.000 348.580 4.300 ;
        RECT 349.740 4.000 350.260 4.300 ;
        RECT 351.420 4.000 351.940 4.300 ;
        RECT 353.100 4.000 353.620 4.300 ;
        RECT 354.780 4.000 355.300 4.300 ;
        RECT 356.460 4.000 356.980 4.300 ;
        RECT 358.140 4.000 358.660 4.300 ;
        RECT 359.820 4.000 360.340 4.300 ;
        RECT 361.500 4.000 362.020 4.300 ;
        RECT 363.180 4.000 363.700 4.300 ;
        RECT 364.860 4.000 365.380 4.300 ;
        RECT 366.540 4.000 367.060 4.300 ;
        RECT 368.220 4.000 368.740 4.300 ;
        RECT 369.900 4.000 370.420 4.300 ;
        RECT 371.580 4.000 372.100 4.300 ;
        RECT 373.260 4.000 373.780 4.300 ;
        RECT 374.940 4.000 375.460 4.300 ;
        RECT 376.620 4.000 377.140 4.300 ;
        RECT 378.300 4.000 378.820 4.300 ;
        RECT 379.980 4.000 380.500 4.300 ;
        RECT 381.660 4.000 382.180 4.300 ;
        RECT 383.340 4.000 383.860 4.300 ;
        RECT 385.020 4.000 385.540 4.300 ;
        RECT 386.700 4.000 387.220 4.300 ;
        RECT 388.380 4.000 388.900 4.300 ;
        RECT 390.060 4.000 390.580 4.300 ;
        RECT 391.740 4.000 392.260 4.300 ;
        RECT 393.420 4.000 393.940 4.300 ;
        RECT 395.100 4.000 395.620 4.300 ;
        RECT 396.780 4.000 397.300 4.300 ;
        RECT 398.460 4.000 398.980 4.300 ;
        RECT 400.140 4.000 400.660 4.300 ;
        RECT 401.820 4.000 402.340 4.300 ;
        RECT 403.500 4.000 404.020 4.300 ;
        RECT 405.180 4.000 405.700 4.300 ;
        RECT 406.860 4.000 407.380 4.300 ;
        RECT 408.540 4.000 409.060 4.300 ;
        RECT 410.220 4.000 410.740 4.300 ;
        RECT 411.900 4.000 412.420 4.300 ;
        RECT 413.580 4.000 414.100 4.300 ;
        RECT 415.260 4.000 415.780 4.300 ;
        RECT 416.940 4.000 417.460 4.300 ;
        RECT 418.620 4.000 419.140 4.300 ;
        RECT 420.300 4.000 420.820 4.300 ;
        RECT 421.980 4.000 422.500 4.300 ;
        RECT 423.660 4.000 424.180 4.300 ;
        RECT 425.340 4.000 425.860 4.300 ;
        RECT 427.020 4.000 427.540 4.300 ;
        RECT 428.700 4.000 429.220 4.300 ;
        RECT 430.380 4.000 430.900 4.300 ;
        RECT 432.060 4.000 432.580 4.300 ;
        RECT 433.740 4.000 434.260 4.300 ;
        RECT 435.420 4.000 435.940 4.300 ;
        RECT 437.100 4.000 437.620 4.300 ;
        RECT 438.780 4.000 439.300 4.300 ;
        RECT 440.460 4.000 440.980 4.300 ;
        RECT 442.140 4.000 442.660 4.300 ;
        RECT 443.820 4.000 444.340 4.300 ;
        RECT 445.500 4.000 446.020 4.300 ;
        RECT 447.180 4.000 447.700 4.300 ;
        RECT 448.860 4.000 449.380 4.300 ;
        RECT 450.540 4.000 451.060 4.300 ;
        RECT 452.220 4.000 452.740 4.300 ;
        RECT 453.900 4.000 454.420 4.300 ;
        RECT 455.580 4.000 456.100 4.300 ;
        RECT 457.260 4.000 457.780 4.300 ;
        RECT 458.940 4.000 459.460 4.300 ;
        RECT 460.620 4.000 461.140 4.300 ;
        RECT 462.300 4.000 462.820 4.300 ;
        RECT 463.980 4.000 464.500 4.300 ;
        RECT 465.660 4.000 466.180 4.300 ;
        RECT 467.340 4.000 467.860 4.300 ;
        RECT 469.020 4.000 469.540 4.300 ;
        RECT 470.700 4.000 471.220 4.300 ;
        RECT 472.380 4.000 472.900 4.300 ;
        RECT 474.060 4.000 474.580 4.300 ;
        RECT 475.740 4.000 476.260 4.300 ;
        RECT 477.420 4.000 477.940 4.300 ;
        RECT 479.100 4.000 479.620 4.300 ;
        RECT 480.780 4.000 481.300 4.300 ;
        RECT 482.460 4.000 482.980 4.300 ;
        RECT 484.140 4.000 484.660 4.300 ;
        RECT 485.820 4.000 486.340 4.300 ;
        RECT 487.500 4.000 488.020 4.300 ;
        RECT 489.180 4.000 489.700 4.300 ;
        RECT 490.860 4.000 491.380 4.300 ;
        RECT 492.540 4.000 493.060 4.300 ;
        RECT 494.220 4.000 494.740 4.300 ;
        RECT 495.900 4.000 496.420 4.300 ;
        RECT 497.580 4.000 498.100 4.300 ;
        RECT 499.260 4.000 499.780 4.300 ;
        RECT 500.940 4.000 501.460 4.300 ;
        RECT 502.620 4.000 503.140 4.300 ;
        RECT 504.300 4.000 504.820 4.300 ;
        RECT 505.980 4.000 506.500 4.300 ;
        RECT 507.660 4.000 508.180 4.300 ;
        RECT 509.340 4.000 509.860 4.300 ;
        RECT 511.020 4.000 511.540 4.300 ;
        RECT 512.700 4.000 513.220 4.300 ;
        RECT 514.380 4.000 514.900 4.300 ;
        RECT 516.060 4.000 516.580 4.300 ;
        RECT 517.740 4.000 518.260 4.300 ;
        RECT 519.420 4.000 519.940 4.300 ;
        RECT 521.100 4.000 521.620 4.300 ;
        RECT 522.780 4.000 523.300 4.300 ;
        RECT 524.460 4.000 524.980 4.300 ;
        RECT 526.140 4.000 526.660 4.300 ;
        RECT 527.820 4.000 528.340 4.300 ;
        RECT 529.500 4.000 530.020 4.300 ;
        RECT 531.180 4.000 531.700 4.300 ;
        RECT 532.860 4.000 533.380 4.300 ;
        RECT 534.540 4.000 535.060 4.300 ;
        RECT 536.220 4.000 536.740 4.300 ;
        RECT 537.900 4.000 538.420 4.300 ;
        RECT 539.580 4.000 540.100 4.300 ;
        RECT 541.260 4.000 541.780 4.300 ;
        RECT 542.940 4.000 543.460 4.300 ;
        RECT 544.620 4.000 545.140 4.300 ;
        RECT 546.300 4.000 546.820 4.300 ;
        RECT 547.980 4.000 548.500 4.300 ;
        RECT 549.660 4.000 588.420 4.300 ;
      LAYER Metal3 ;
        RECT 20.810 8.540 577.830 588.420 ;
      LAYER Metal4 ;
        RECT 226.380 551.130 252.340 582.310 ;
        RECT 254.540 551.130 329.140 582.310 ;
        RECT 331.340 551.130 394.660 582.310 ;
  END
END macro_golden
END LIBRARY

