magic
tech gf180mcuC
magscale 1 5
timestamp 1670058194
<< obsm1 >>
rect 672 855 89320 58785
<< metal2 >>
rect 3472 59600 3528 60000
rect 4200 59600 4256 60000
rect 4928 59600 4984 60000
rect 5656 59600 5712 60000
rect 6384 59600 6440 60000
rect 7112 59600 7168 60000
rect 7840 59600 7896 60000
rect 8568 59600 8624 60000
rect 9296 59600 9352 60000
rect 10024 59600 10080 60000
rect 10752 59600 10808 60000
rect 11480 59600 11536 60000
rect 12208 59600 12264 60000
rect 12936 59600 12992 60000
rect 13664 59600 13720 60000
rect 14392 59600 14448 60000
rect 15120 59600 15176 60000
rect 15848 59600 15904 60000
rect 16576 59600 16632 60000
rect 17304 59600 17360 60000
rect 18032 59600 18088 60000
rect 18760 59600 18816 60000
rect 19488 59600 19544 60000
rect 20216 59600 20272 60000
rect 20944 59600 21000 60000
rect 21672 59600 21728 60000
rect 22400 59600 22456 60000
rect 23128 59600 23184 60000
rect 23856 59600 23912 60000
rect 24584 59600 24640 60000
rect 25312 59600 25368 60000
rect 26040 59600 26096 60000
rect 26768 59600 26824 60000
rect 27496 59600 27552 60000
rect 28224 59600 28280 60000
rect 28952 59600 29008 60000
rect 29680 59600 29736 60000
rect 30408 59600 30464 60000
rect 31136 59600 31192 60000
rect 31864 59600 31920 60000
rect 32592 59600 32648 60000
rect 33320 59600 33376 60000
rect 34048 59600 34104 60000
rect 34776 59600 34832 60000
rect 35504 59600 35560 60000
rect 36232 59600 36288 60000
rect 36960 59600 37016 60000
rect 37688 59600 37744 60000
rect 38416 59600 38472 60000
rect 39144 59600 39200 60000
rect 39872 59600 39928 60000
rect 40600 59600 40656 60000
rect 41328 59600 41384 60000
rect 42056 59600 42112 60000
rect 42784 59600 42840 60000
rect 43512 59600 43568 60000
rect 44240 59600 44296 60000
rect 44968 59600 45024 60000
rect 45696 59600 45752 60000
rect 46424 59600 46480 60000
rect 47152 59600 47208 60000
rect 47880 59600 47936 60000
rect 48608 59600 48664 60000
rect 49336 59600 49392 60000
rect 50064 59600 50120 60000
rect 50792 59600 50848 60000
rect 51520 59600 51576 60000
rect 52248 59600 52304 60000
rect 52976 59600 53032 60000
rect 53704 59600 53760 60000
rect 54432 59600 54488 60000
rect 55160 59600 55216 60000
rect 55888 59600 55944 60000
rect 56616 59600 56672 60000
rect 57344 59600 57400 60000
rect 58072 59600 58128 60000
rect 58800 59600 58856 60000
rect 59528 59600 59584 60000
rect 60256 59600 60312 60000
rect 60984 59600 61040 60000
rect 61712 59600 61768 60000
rect 62440 59600 62496 60000
rect 63168 59600 63224 60000
rect 63896 59600 63952 60000
rect 64624 59600 64680 60000
rect 65352 59600 65408 60000
rect 66080 59600 66136 60000
rect 66808 59600 66864 60000
rect 67536 59600 67592 60000
rect 68264 59600 68320 60000
rect 68992 59600 69048 60000
rect 69720 59600 69776 60000
rect 70448 59600 70504 60000
rect 71176 59600 71232 60000
rect 71904 59600 71960 60000
rect 72632 59600 72688 60000
rect 73360 59600 73416 60000
rect 74088 59600 74144 60000
rect 74816 59600 74872 60000
rect 75544 59600 75600 60000
rect 76272 59600 76328 60000
rect 77000 59600 77056 60000
rect 77728 59600 77784 60000
rect 78456 59600 78512 60000
rect 79184 59600 79240 60000
rect 79912 59600 79968 60000
rect 80640 59600 80696 60000
rect 81368 59600 81424 60000
rect 82096 59600 82152 60000
rect 82824 59600 82880 60000
rect 83552 59600 83608 60000
rect 84280 59600 84336 60000
rect 85008 59600 85064 60000
rect 85736 59600 85792 60000
rect 86464 59600 86520 60000
rect 3864 0 3920 400
rect 4032 0 4088 400
rect 4200 0 4256 400
rect 4368 0 4424 400
rect 4536 0 4592 400
rect 4704 0 4760 400
rect 4872 0 4928 400
rect 5040 0 5096 400
rect 5208 0 5264 400
rect 5376 0 5432 400
rect 5544 0 5600 400
rect 5712 0 5768 400
rect 5880 0 5936 400
rect 6048 0 6104 400
rect 6216 0 6272 400
rect 6384 0 6440 400
rect 6552 0 6608 400
rect 6720 0 6776 400
rect 6888 0 6944 400
rect 7056 0 7112 400
rect 7224 0 7280 400
rect 7392 0 7448 400
rect 7560 0 7616 400
rect 7728 0 7784 400
rect 7896 0 7952 400
rect 8064 0 8120 400
rect 8232 0 8288 400
rect 8400 0 8456 400
rect 8568 0 8624 400
rect 8736 0 8792 400
rect 8904 0 8960 400
rect 9072 0 9128 400
rect 9240 0 9296 400
rect 9408 0 9464 400
rect 9576 0 9632 400
rect 9744 0 9800 400
rect 9912 0 9968 400
rect 10080 0 10136 400
rect 10248 0 10304 400
rect 10416 0 10472 400
rect 10584 0 10640 400
rect 10752 0 10808 400
rect 10920 0 10976 400
rect 11088 0 11144 400
rect 11256 0 11312 400
rect 11424 0 11480 400
rect 11592 0 11648 400
rect 11760 0 11816 400
rect 11928 0 11984 400
rect 12096 0 12152 400
rect 12264 0 12320 400
rect 12432 0 12488 400
rect 12600 0 12656 400
rect 12768 0 12824 400
rect 12936 0 12992 400
rect 13104 0 13160 400
rect 13272 0 13328 400
rect 13440 0 13496 400
rect 13608 0 13664 400
rect 13776 0 13832 400
rect 13944 0 14000 400
rect 14112 0 14168 400
rect 14280 0 14336 400
rect 14448 0 14504 400
rect 14616 0 14672 400
rect 14784 0 14840 400
rect 14952 0 15008 400
rect 15120 0 15176 400
rect 15288 0 15344 400
rect 15456 0 15512 400
rect 15624 0 15680 400
rect 15792 0 15848 400
rect 15960 0 16016 400
rect 16128 0 16184 400
rect 16296 0 16352 400
rect 16464 0 16520 400
rect 16632 0 16688 400
rect 16800 0 16856 400
rect 16968 0 17024 400
rect 17136 0 17192 400
rect 17304 0 17360 400
rect 17472 0 17528 400
rect 17640 0 17696 400
rect 17808 0 17864 400
rect 17976 0 18032 400
rect 18144 0 18200 400
rect 18312 0 18368 400
rect 18480 0 18536 400
rect 18648 0 18704 400
rect 18816 0 18872 400
rect 18984 0 19040 400
rect 19152 0 19208 400
rect 19320 0 19376 400
rect 19488 0 19544 400
rect 19656 0 19712 400
rect 19824 0 19880 400
rect 19992 0 20048 400
rect 20160 0 20216 400
rect 20328 0 20384 400
rect 20496 0 20552 400
rect 20664 0 20720 400
rect 20832 0 20888 400
rect 21000 0 21056 400
rect 21168 0 21224 400
rect 21336 0 21392 400
rect 21504 0 21560 400
rect 21672 0 21728 400
rect 21840 0 21896 400
rect 22008 0 22064 400
rect 22176 0 22232 400
rect 22344 0 22400 400
rect 22512 0 22568 400
rect 22680 0 22736 400
rect 22848 0 22904 400
rect 23016 0 23072 400
rect 23184 0 23240 400
rect 23352 0 23408 400
rect 23520 0 23576 400
rect 23688 0 23744 400
rect 23856 0 23912 400
rect 24024 0 24080 400
rect 24192 0 24248 400
rect 24360 0 24416 400
rect 24528 0 24584 400
rect 24696 0 24752 400
rect 24864 0 24920 400
rect 25032 0 25088 400
rect 25200 0 25256 400
rect 25368 0 25424 400
rect 25536 0 25592 400
rect 25704 0 25760 400
rect 25872 0 25928 400
rect 26040 0 26096 400
rect 26208 0 26264 400
rect 26376 0 26432 400
rect 26544 0 26600 400
rect 26712 0 26768 400
rect 26880 0 26936 400
rect 27048 0 27104 400
rect 27216 0 27272 400
rect 27384 0 27440 400
rect 27552 0 27608 400
rect 27720 0 27776 400
rect 27888 0 27944 400
rect 28056 0 28112 400
rect 28224 0 28280 400
rect 28392 0 28448 400
rect 28560 0 28616 400
rect 28728 0 28784 400
rect 28896 0 28952 400
rect 29064 0 29120 400
rect 29232 0 29288 400
rect 29400 0 29456 400
rect 29568 0 29624 400
rect 29736 0 29792 400
rect 29904 0 29960 400
rect 30072 0 30128 400
rect 30240 0 30296 400
rect 30408 0 30464 400
rect 30576 0 30632 400
rect 30744 0 30800 400
rect 30912 0 30968 400
rect 31080 0 31136 400
rect 31248 0 31304 400
rect 31416 0 31472 400
rect 31584 0 31640 400
rect 31752 0 31808 400
rect 31920 0 31976 400
rect 32088 0 32144 400
rect 32256 0 32312 400
rect 32424 0 32480 400
rect 32592 0 32648 400
rect 32760 0 32816 400
rect 32928 0 32984 400
rect 33096 0 33152 400
rect 33264 0 33320 400
rect 33432 0 33488 400
rect 33600 0 33656 400
rect 33768 0 33824 400
rect 33936 0 33992 400
rect 34104 0 34160 400
rect 34272 0 34328 400
rect 34440 0 34496 400
rect 34608 0 34664 400
rect 34776 0 34832 400
rect 34944 0 35000 400
rect 35112 0 35168 400
rect 35280 0 35336 400
rect 35448 0 35504 400
rect 35616 0 35672 400
rect 35784 0 35840 400
rect 35952 0 36008 400
rect 36120 0 36176 400
rect 36288 0 36344 400
rect 36456 0 36512 400
rect 36624 0 36680 400
rect 36792 0 36848 400
rect 36960 0 37016 400
rect 37128 0 37184 400
rect 37296 0 37352 400
rect 37464 0 37520 400
rect 37632 0 37688 400
rect 37800 0 37856 400
rect 37968 0 38024 400
rect 38136 0 38192 400
rect 38304 0 38360 400
rect 38472 0 38528 400
rect 38640 0 38696 400
rect 38808 0 38864 400
rect 38976 0 39032 400
rect 39144 0 39200 400
rect 39312 0 39368 400
rect 39480 0 39536 400
rect 39648 0 39704 400
rect 39816 0 39872 400
rect 39984 0 40040 400
rect 40152 0 40208 400
rect 40320 0 40376 400
rect 40488 0 40544 400
rect 40656 0 40712 400
rect 40824 0 40880 400
rect 40992 0 41048 400
rect 41160 0 41216 400
rect 41328 0 41384 400
rect 41496 0 41552 400
rect 41664 0 41720 400
rect 41832 0 41888 400
rect 42000 0 42056 400
rect 42168 0 42224 400
rect 42336 0 42392 400
rect 42504 0 42560 400
rect 42672 0 42728 400
rect 42840 0 42896 400
rect 43008 0 43064 400
rect 43176 0 43232 400
rect 43344 0 43400 400
rect 43512 0 43568 400
rect 43680 0 43736 400
rect 43848 0 43904 400
rect 44016 0 44072 400
rect 44184 0 44240 400
rect 44352 0 44408 400
rect 44520 0 44576 400
rect 44688 0 44744 400
rect 44856 0 44912 400
rect 45024 0 45080 400
rect 45192 0 45248 400
rect 45360 0 45416 400
rect 45528 0 45584 400
rect 45696 0 45752 400
rect 45864 0 45920 400
rect 46032 0 46088 400
rect 46200 0 46256 400
rect 46368 0 46424 400
rect 46536 0 46592 400
rect 46704 0 46760 400
rect 46872 0 46928 400
rect 47040 0 47096 400
rect 47208 0 47264 400
rect 47376 0 47432 400
rect 47544 0 47600 400
rect 47712 0 47768 400
rect 47880 0 47936 400
rect 48048 0 48104 400
rect 48216 0 48272 400
rect 48384 0 48440 400
rect 48552 0 48608 400
rect 48720 0 48776 400
rect 48888 0 48944 400
rect 49056 0 49112 400
rect 49224 0 49280 400
rect 49392 0 49448 400
rect 49560 0 49616 400
rect 49728 0 49784 400
rect 49896 0 49952 400
rect 50064 0 50120 400
rect 50232 0 50288 400
rect 50400 0 50456 400
rect 50568 0 50624 400
rect 50736 0 50792 400
rect 50904 0 50960 400
rect 51072 0 51128 400
rect 51240 0 51296 400
rect 51408 0 51464 400
rect 51576 0 51632 400
rect 51744 0 51800 400
rect 51912 0 51968 400
rect 52080 0 52136 400
rect 52248 0 52304 400
rect 52416 0 52472 400
rect 52584 0 52640 400
rect 52752 0 52808 400
rect 52920 0 52976 400
rect 53088 0 53144 400
rect 53256 0 53312 400
rect 53424 0 53480 400
rect 53592 0 53648 400
rect 53760 0 53816 400
rect 53928 0 53984 400
rect 54096 0 54152 400
rect 54264 0 54320 400
rect 54432 0 54488 400
rect 54600 0 54656 400
rect 54768 0 54824 400
rect 54936 0 54992 400
rect 55104 0 55160 400
rect 55272 0 55328 400
rect 55440 0 55496 400
rect 55608 0 55664 400
rect 55776 0 55832 400
rect 55944 0 56000 400
rect 56112 0 56168 400
rect 56280 0 56336 400
rect 56448 0 56504 400
rect 56616 0 56672 400
rect 56784 0 56840 400
rect 56952 0 57008 400
rect 57120 0 57176 400
rect 57288 0 57344 400
rect 57456 0 57512 400
rect 57624 0 57680 400
rect 57792 0 57848 400
rect 57960 0 58016 400
rect 58128 0 58184 400
rect 58296 0 58352 400
rect 58464 0 58520 400
rect 58632 0 58688 400
rect 58800 0 58856 400
rect 58968 0 59024 400
rect 59136 0 59192 400
rect 59304 0 59360 400
rect 59472 0 59528 400
rect 59640 0 59696 400
rect 59808 0 59864 400
rect 59976 0 60032 400
rect 60144 0 60200 400
rect 60312 0 60368 400
rect 60480 0 60536 400
rect 60648 0 60704 400
rect 60816 0 60872 400
rect 60984 0 61040 400
rect 61152 0 61208 400
rect 61320 0 61376 400
rect 61488 0 61544 400
rect 61656 0 61712 400
rect 61824 0 61880 400
rect 61992 0 62048 400
rect 62160 0 62216 400
rect 62328 0 62384 400
rect 62496 0 62552 400
rect 62664 0 62720 400
rect 62832 0 62888 400
rect 63000 0 63056 400
rect 63168 0 63224 400
rect 63336 0 63392 400
rect 63504 0 63560 400
rect 63672 0 63728 400
rect 63840 0 63896 400
rect 64008 0 64064 400
rect 64176 0 64232 400
rect 64344 0 64400 400
rect 64512 0 64568 400
rect 64680 0 64736 400
rect 64848 0 64904 400
rect 65016 0 65072 400
rect 65184 0 65240 400
rect 65352 0 65408 400
rect 65520 0 65576 400
rect 65688 0 65744 400
rect 65856 0 65912 400
rect 66024 0 66080 400
rect 66192 0 66248 400
rect 66360 0 66416 400
rect 66528 0 66584 400
rect 66696 0 66752 400
rect 66864 0 66920 400
rect 67032 0 67088 400
rect 67200 0 67256 400
rect 67368 0 67424 400
rect 67536 0 67592 400
rect 67704 0 67760 400
rect 67872 0 67928 400
rect 68040 0 68096 400
rect 68208 0 68264 400
rect 68376 0 68432 400
rect 68544 0 68600 400
rect 68712 0 68768 400
rect 68880 0 68936 400
rect 69048 0 69104 400
rect 69216 0 69272 400
rect 69384 0 69440 400
rect 69552 0 69608 400
rect 69720 0 69776 400
rect 69888 0 69944 400
rect 70056 0 70112 400
rect 70224 0 70280 400
rect 70392 0 70448 400
rect 70560 0 70616 400
rect 70728 0 70784 400
rect 70896 0 70952 400
rect 71064 0 71120 400
rect 71232 0 71288 400
rect 71400 0 71456 400
rect 71568 0 71624 400
rect 71736 0 71792 400
rect 71904 0 71960 400
rect 72072 0 72128 400
rect 72240 0 72296 400
rect 72408 0 72464 400
rect 72576 0 72632 400
rect 72744 0 72800 400
rect 72912 0 72968 400
rect 73080 0 73136 400
rect 73248 0 73304 400
rect 73416 0 73472 400
rect 73584 0 73640 400
rect 73752 0 73808 400
rect 73920 0 73976 400
rect 74088 0 74144 400
rect 74256 0 74312 400
rect 74424 0 74480 400
rect 74592 0 74648 400
rect 74760 0 74816 400
rect 74928 0 74984 400
rect 75096 0 75152 400
rect 75264 0 75320 400
rect 75432 0 75488 400
rect 75600 0 75656 400
rect 75768 0 75824 400
rect 75936 0 75992 400
rect 76104 0 76160 400
rect 76272 0 76328 400
rect 76440 0 76496 400
rect 76608 0 76664 400
rect 76776 0 76832 400
rect 76944 0 77000 400
rect 77112 0 77168 400
rect 77280 0 77336 400
rect 77448 0 77504 400
rect 77616 0 77672 400
rect 77784 0 77840 400
rect 77952 0 78008 400
rect 78120 0 78176 400
rect 78288 0 78344 400
rect 78456 0 78512 400
rect 78624 0 78680 400
rect 78792 0 78848 400
rect 78960 0 79016 400
rect 79128 0 79184 400
rect 79296 0 79352 400
rect 79464 0 79520 400
rect 79632 0 79688 400
rect 79800 0 79856 400
rect 79968 0 80024 400
rect 80136 0 80192 400
rect 80304 0 80360 400
rect 80472 0 80528 400
rect 80640 0 80696 400
rect 80808 0 80864 400
rect 80976 0 81032 400
rect 81144 0 81200 400
rect 81312 0 81368 400
rect 81480 0 81536 400
rect 81648 0 81704 400
rect 81816 0 81872 400
rect 81984 0 82040 400
rect 82152 0 82208 400
rect 82320 0 82376 400
rect 82488 0 82544 400
rect 82656 0 82712 400
rect 82824 0 82880 400
rect 82992 0 83048 400
rect 83160 0 83216 400
rect 83328 0 83384 400
rect 83496 0 83552 400
rect 83664 0 83720 400
rect 83832 0 83888 400
rect 84000 0 84056 400
rect 84168 0 84224 400
rect 84336 0 84392 400
rect 84504 0 84560 400
rect 84672 0 84728 400
rect 84840 0 84896 400
rect 85008 0 85064 400
rect 85176 0 85232 400
rect 85344 0 85400 400
rect 85512 0 85568 400
rect 85680 0 85736 400
rect 85848 0 85904 400
rect 86016 0 86072 400
<< obsm2 >>
rect 2238 59570 3442 59600
rect 3558 59570 4170 59600
rect 4286 59570 4898 59600
rect 5014 59570 5626 59600
rect 5742 59570 6354 59600
rect 6470 59570 7082 59600
rect 7198 59570 7810 59600
rect 7926 59570 8538 59600
rect 8654 59570 9266 59600
rect 9382 59570 9994 59600
rect 10110 59570 10722 59600
rect 10838 59570 11450 59600
rect 11566 59570 12178 59600
rect 12294 59570 12906 59600
rect 13022 59570 13634 59600
rect 13750 59570 14362 59600
rect 14478 59570 15090 59600
rect 15206 59570 15818 59600
rect 15934 59570 16546 59600
rect 16662 59570 17274 59600
rect 17390 59570 18002 59600
rect 18118 59570 18730 59600
rect 18846 59570 19458 59600
rect 19574 59570 20186 59600
rect 20302 59570 20914 59600
rect 21030 59570 21642 59600
rect 21758 59570 22370 59600
rect 22486 59570 23098 59600
rect 23214 59570 23826 59600
rect 23942 59570 24554 59600
rect 24670 59570 25282 59600
rect 25398 59570 26010 59600
rect 26126 59570 26738 59600
rect 26854 59570 27466 59600
rect 27582 59570 28194 59600
rect 28310 59570 28922 59600
rect 29038 59570 29650 59600
rect 29766 59570 30378 59600
rect 30494 59570 31106 59600
rect 31222 59570 31834 59600
rect 31950 59570 32562 59600
rect 32678 59570 33290 59600
rect 33406 59570 34018 59600
rect 34134 59570 34746 59600
rect 34862 59570 35474 59600
rect 35590 59570 36202 59600
rect 36318 59570 36930 59600
rect 37046 59570 37658 59600
rect 37774 59570 38386 59600
rect 38502 59570 39114 59600
rect 39230 59570 39842 59600
rect 39958 59570 40570 59600
rect 40686 59570 41298 59600
rect 41414 59570 42026 59600
rect 42142 59570 42754 59600
rect 42870 59570 43482 59600
rect 43598 59570 44210 59600
rect 44326 59570 44938 59600
rect 45054 59570 45666 59600
rect 45782 59570 46394 59600
rect 46510 59570 47122 59600
rect 47238 59570 47850 59600
rect 47966 59570 48578 59600
rect 48694 59570 49306 59600
rect 49422 59570 50034 59600
rect 50150 59570 50762 59600
rect 50878 59570 51490 59600
rect 51606 59570 52218 59600
rect 52334 59570 52946 59600
rect 53062 59570 53674 59600
rect 53790 59570 54402 59600
rect 54518 59570 55130 59600
rect 55246 59570 55858 59600
rect 55974 59570 56586 59600
rect 56702 59570 57314 59600
rect 57430 59570 58042 59600
rect 58158 59570 58770 59600
rect 58886 59570 59498 59600
rect 59614 59570 60226 59600
rect 60342 59570 60954 59600
rect 61070 59570 61682 59600
rect 61798 59570 62410 59600
rect 62526 59570 63138 59600
rect 63254 59570 63866 59600
rect 63982 59570 64594 59600
rect 64710 59570 65322 59600
rect 65438 59570 66050 59600
rect 66166 59570 66778 59600
rect 66894 59570 67506 59600
rect 67622 59570 68234 59600
rect 68350 59570 68962 59600
rect 69078 59570 69690 59600
rect 69806 59570 70418 59600
rect 70534 59570 71146 59600
rect 71262 59570 71874 59600
rect 71990 59570 72602 59600
rect 72718 59570 73330 59600
rect 73446 59570 74058 59600
rect 74174 59570 74786 59600
rect 74902 59570 75514 59600
rect 75630 59570 76242 59600
rect 76358 59570 76970 59600
rect 77086 59570 77698 59600
rect 77814 59570 78426 59600
rect 78542 59570 79154 59600
rect 79270 59570 79882 59600
rect 79998 59570 80610 59600
rect 80726 59570 81338 59600
rect 81454 59570 82066 59600
rect 82182 59570 82794 59600
rect 82910 59570 83522 59600
rect 83638 59570 84250 59600
rect 84366 59570 84978 59600
rect 85094 59570 85706 59600
rect 85822 59570 86434 59600
rect 86550 59570 86850 59600
rect 2238 430 86850 59570
rect 2238 400 3834 430
rect 3950 400 4002 430
rect 4118 400 4170 430
rect 4286 400 4338 430
rect 4454 400 4506 430
rect 4622 400 4674 430
rect 4790 400 4842 430
rect 4958 400 5010 430
rect 5126 400 5178 430
rect 5294 400 5346 430
rect 5462 400 5514 430
rect 5630 400 5682 430
rect 5798 400 5850 430
rect 5966 400 6018 430
rect 6134 400 6186 430
rect 6302 400 6354 430
rect 6470 400 6522 430
rect 6638 400 6690 430
rect 6806 400 6858 430
rect 6974 400 7026 430
rect 7142 400 7194 430
rect 7310 400 7362 430
rect 7478 400 7530 430
rect 7646 400 7698 430
rect 7814 400 7866 430
rect 7982 400 8034 430
rect 8150 400 8202 430
rect 8318 400 8370 430
rect 8486 400 8538 430
rect 8654 400 8706 430
rect 8822 400 8874 430
rect 8990 400 9042 430
rect 9158 400 9210 430
rect 9326 400 9378 430
rect 9494 400 9546 430
rect 9662 400 9714 430
rect 9830 400 9882 430
rect 9998 400 10050 430
rect 10166 400 10218 430
rect 10334 400 10386 430
rect 10502 400 10554 430
rect 10670 400 10722 430
rect 10838 400 10890 430
rect 11006 400 11058 430
rect 11174 400 11226 430
rect 11342 400 11394 430
rect 11510 400 11562 430
rect 11678 400 11730 430
rect 11846 400 11898 430
rect 12014 400 12066 430
rect 12182 400 12234 430
rect 12350 400 12402 430
rect 12518 400 12570 430
rect 12686 400 12738 430
rect 12854 400 12906 430
rect 13022 400 13074 430
rect 13190 400 13242 430
rect 13358 400 13410 430
rect 13526 400 13578 430
rect 13694 400 13746 430
rect 13862 400 13914 430
rect 14030 400 14082 430
rect 14198 400 14250 430
rect 14366 400 14418 430
rect 14534 400 14586 430
rect 14702 400 14754 430
rect 14870 400 14922 430
rect 15038 400 15090 430
rect 15206 400 15258 430
rect 15374 400 15426 430
rect 15542 400 15594 430
rect 15710 400 15762 430
rect 15878 400 15930 430
rect 16046 400 16098 430
rect 16214 400 16266 430
rect 16382 400 16434 430
rect 16550 400 16602 430
rect 16718 400 16770 430
rect 16886 400 16938 430
rect 17054 400 17106 430
rect 17222 400 17274 430
rect 17390 400 17442 430
rect 17558 400 17610 430
rect 17726 400 17778 430
rect 17894 400 17946 430
rect 18062 400 18114 430
rect 18230 400 18282 430
rect 18398 400 18450 430
rect 18566 400 18618 430
rect 18734 400 18786 430
rect 18902 400 18954 430
rect 19070 400 19122 430
rect 19238 400 19290 430
rect 19406 400 19458 430
rect 19574 400 19626 430
rect 19742 400 19794 430
rect 19910 400 19962 430
rect 20078 400 20130 430
rect 20246 400 20298 430
rect 20414 400 20466 430
rect 20582 400 20634 430
rect 20750 400 20802 430
rect 20918 400 20970 430
rect 21086 400 21138 430
rect 21254 400 21306 430
rect 21422 400 21474 430
rect 21590 400 21642 430
rect 21758 400 21810 430
rect 21926 400 21978 430
rect 22094 400 22146 430
rect 22262 400 22314 430
rect 22430 400 22482 430
rect 22598 400 22650 430
rect 22766 400 22818 430
rect 22934 400 22986 430
rect 23102 400 23154 430
rect 23270 400 23322 430
rect 23438 400 23490 430
rect 23606 400 23658 430
rect 23774 400 23826 430
rect 23942 400 23994 430
rect 24110 400 24162 430
rect 24278 400 24330 430
rect 24446 400 24498 430
rect 24614 400 24666 430
rect 24782 400 24834 430
rect 24950 400 25002 430
rect 25118 400 25170 430
rect 25286 400 25338 430
rect 25454 400 25506 430
rect 25622 400 25674 430
rect 25790 400 25842 430
rect 25958 400 26010 430
rect 26126 400 26178 430
rect 26294 400 26346 430
rect 26462 400 26514 430
rect 26630 400 26682 430
rect 26798 400 26850 430
rect 26966 400 27018 430
rect 27134 400 27186 430
rect 27302 400 27354 430
rect 27470 400 27522 430
rect 27638 400 27690 430
rect 27806 400 27858 430
rect 27974 400 28026 430
rect 28142 400 28194 430
rect 28310 400 28362 430
rect 28478 400 28530 430
rect 28646 400 28698 430
rect 28814 400 28866 430
rect 28982 400 29034 430
rect 29150 400 29202 430
rect 29318 400 29370 430
rect 29486 400 29538 430
rect 29654 400 29706 430
rect 29822 400 29874 430
rect 29990 400 30042 430
rect 30158 400 30210 430
rect 30326 400 30378 430
rect 30494 400 30546 430
rect 30662 400 30714 430
rect 30830 400 30882 430
rect 30998 400 31050 430
rect 31166 400 31218 430
rect 31334 400 31386 430
rect 31502 400 31554 430
rect 31670 400 31722 430
rect 31838 400 31890 430
rect 32006 400 32058 430
rect 32174 400 32226 430
rect 32342 400 32394 430
rect 32510 400 32562 430
rect 32678 400 32730 430
rect 32846 400 32898 430
rect 33014 400 33066 430
rect 33182 400 33234 430
rect 33350 400 33402 430
rect 33518 400 33570 430
rect 33686 400 33738 430
rect 33854 400 33906 430
rect 34022 400 34074 430
rect 34190 400 34242 430
rect 34358 400 34410 430
rect 34526 400 34578 430
rect 34694 400 34746 430
rect 34862 400 34914 430
rect 35030 400 35082 430
rect 35198 400 35250 430
rect 35366 400 35418 430
rect 35534 400 35586 430
rect 35702 400 35754 430
rect 35870 400 35922 430
rect 36038 400 36090 430
rect 36206 400 36258 430
rect 36374 400 36426 430
rect 36542 400 36594 430
rect 36710 400 36762 430
rect 36878 400 36930 430
rect 37046 400 37098 430
rect 37214 400 37266 430
rect 37382 400 37434 430
rect 37550 400 37602 430
rect 37718 400 37770 430
rect 37886 400 37938 430
rect 38054 400 38106 430
rect 38222 400 38274 430
rect 38390 400 38442 430
rect 38558 400 38610 430
rect 38726 400 38778 430
rect 38894 400 38946 430
rect 39062 400 39114 430
rect 39230 400 39282 430
rect 39398 400 39450 430
rect 39566 400 39618 430
rect 39734 400 39786 430
rect 39902 400 39954 430
rect 40070 400 40122 430
rect 40238 400 40290 430
rect 40406 400 40458 430
rect 40574 400 40626 430
rect 40742 400 40794 430
rect 40910 400 40962 430
rect 41078 400 41130 430
rect 41246 400 41298 430
rect 41414 400 41466 430
rect 41582 400 41634 430
rect 41750 400 41802 430
rect 41918 400 41970 430
rect 42086 400 42138 430
rect 42254 400 42306 430
rect 42422 400 42474 430
rect 42590 400 42642 430
rect 42758 400 42810 430
rect 42926 400 42978 430
rect 43094 400 43146 430
rect 43262 400 43314 430
rect 43430 400 43482 430
rect 43598 400 43650 430
rect 43766 400 43818 430
rect 43934 400 43986 430
rect 44102 400 44154 430
rect 44270 400 44322 430
rect 44438 400 44490 430
rect 44606 400 44658 430
rect 44774 400 44826 430
rect 44942 400 44994 430
rect 45110 400 45162 430
rect 45278 400 45330 430
rect 45446 400 45498 430
rect 45614 400 45666 430
rect 45782 400 45834 430
rect 45950 400 46002 430
rect 46118 400 46170 430
rect 46286 400 46338 430
rect 46454 400 46506 430
rect 46622 400 46674 430
rect 46790 400 46842 430
rect 46958 400 47010 430
rect 47126 400 47178 430
rect 47294 400 47346 430
rect 47462 400 47514 430
rect 47630 400 47682 430
rect 47798 400 47850 430
rect 47966 400 48018 430
rect 48134 400 48186 430
rect 48302 400 48354 430
rect 48470 400 48522 430
rect 48638 400 48690 430
rect 48806 400 48858 430
rect 48974 400 49026 430
rect 49142 400 49194 430
rect 49310 400 49362 430
rect 49478 400 49530 430
rect 49646 400 49698 430
rect 49814 400 49866 430
rect 49982 400 50034 430
rect 50150 400 50202 430
rect 50318 400 50370 430
rect 50486 400 50538 430
rect 50654 400 50706 430
rect 50822 400 50874 430
rect 50990 400 51042 430
rect 51158 400 51210 430
rect 51326 400 51378 430
rect 51494 400 51546 430
rect 51662 400 51714 430
rect 51830 400 51882 430
rect 51998 400 52050 430
rect 52166 400 52218 430
rect 52334 400 52386 430
rect 52502 400 52554 430
rect 52670 400 52722 430
rect 52838 400 52890 430
rect 53006 400 53058 430
rect 53174 400 53226 430
rect 53342 400 53394 430
rect 53510 400 53562 430
rect 53678 400 53730 430
rect 53846 400 53898 430
rect 54014 400 54066 430
rect 54182 400 54234 430
rect 54350 400 54402 430
rect 54518 400 54570 430
rect 54686 400 54738 430
rect 54854 400 54906 430
rect 55022 400 55074 430
rect 55190 400 55242 430
rect 55358 400 55410 430
rect 55526 400 55578 430
rect 55694 400 55746 430
rect 55862 400 55914 430
rect 56030 400 56082 430
rect 56198 400 56250 430
rect 56366 400 56418 430
rect 56534 400 56586 430
rect 56702 400 56754 430
rect 56870 400 56922 430
rect 57038 400 57090 430
rect 57206 400 57258 430
rect 57374 400 57426 430
rect 57542 400 57594 430
rect 57710 400 57762 430
rect 57878 400 57930 430
rect 58046 400 58098 430
rect 58214 400 58266 430
rect 58382 400 58434 430
rect 58550 400 58602 430
rect 58718 400 58770 430
rect 58886 400 58938 430
rect 59054 400 59106 430
rect 59222 400 59274 430
rect 59390 400 59442 430
rect 59558 400 59610 430
rect 59726 400 59778 430
rect 59894 400 59946 430
rect 60062 400 60114 430
rect 60230 400 60282 430
rect 60398 400 60450 430
rect 60566 400 60618 430
rect 60734 400 60786 430
rect 60902 400 60954 430
rect 61070 400 61122 430
rect 61238 400 61290 430
rect 61406 400 61458 430
rect 61574 400 61626 430
rect 61742 400 61794 430
rect 61910 400 61962 430
rect 62078 400 62130 430
rect 62246 400 62298 430
rect 62414 400 62466 430
rect 62582 400 62634 430
rect 62750 400 62802 430
rect 62918 400 62970 430
rect 63086 400 63138 430
rect 63254 400 63306 430
rect 63422 400 63474 430
rect 63590 400 63642 430
rect 63758 400 63810 430
rect 63926 400 63978 430
rect 64094 400 64146 430
rect 64262 400 64314 430
rect 64430 400 64482 430
rect 64598 400 64650 430
rect 64766 400 64818 430
rect 64934 400 64986 430
rect 65102 400 65154 430
rect 65270 400 65322 430
rect 65438 400 65490 430
rect 65606 400 65658 430
rect 65774 400 65826 430
rect 65942 400 65994 430
rect 66110 400 66162 430
rect 66278 400 66330 430
rect 66446 400 66498 430
rect 66614 400 66666 430
rect 66782 400 66834 430
rect 66950 400 67002 430
rect 67118 400 67170 430
rect 67286 400 67338 430
rect 67454 400 67506 430
rect 67622 400 67674 430
rect 67790 400 67842 430
rect 67958 400 68010 430
rect 68126 400 68178 430
rect 68294 400 68346 430
rect 68462 400 68514 430
rect 68630 400 68682 430
rect 68798 400 68850 430
rect 68966 400 69018 430
rect 69134 400 69186 430
rect 69302 400 69354 430
rect 69470 400 69522 430
rect 69638 400 69690 430
rect 69806 400 69858 430
rect 69974 400 70026 430
rect 70142 400 70194 430
rect 70310 400 70362 430
rect 70478 400 70530 430
rect 70646 400 70698 430
rect 70814 400 70866 430
rect 70982 400 71034 430
rect 71150 400 71202 430
rect 71318 400 71370 430
rect 71486 400 71538 430
rect 71654 400 71706 430
rect 71822 400 71874 430
rect 71990 400 72042 430
rect 72158 400 72210 430
rect 72326 400 72378 430
rect 72494 400 72546 430
rect 72662 400 72714 430
rect 72830 400 72882 430
rect 72998 400 73050 430
rect 73166 400 73218 430
rect 73334 400 73386 430
rect 73502 400 73554 430
rect 73670 400 73722 430
rect 73838 400 73890 430
rect 74006 400 74058 430
rect 74174 400 74226 430
rect 74342 400 74394 430
rect 74510 400 74562 430
rect 74678 400 74730 430
rect 74846 400 74898 430
rect 75014 400 75066 430
rect 75182 400 75234 430
rect 75350 400 75402 430
rect 75518 400 75570 430
rect 75686 400 75738 430
rect 75854 400 75906 430
rect 76022 400 76074 430
rect 76190 400 76242 430
rect 76358 400 76410 430
rect 76526 400 76578 430
rect 76694 400 76746 430
rect 76862 400 76914 430
rect 77030 400 77082 430
rect 77198 400 77250 430
rect 77366 400 77418 430
rect 77534 400 77586 430
rect 77702 400 77754 430
rect 77870 400 77922 430
rect 78038 400 78090 430
rect 78206 400 78258 430
rect 78374 400 78426 430
rect 78542 400 78594 430
rect 78710 400 78762 430
rect 78878 400 78930 430
rect 79046 400 79098 430
rect 79214 400 79266 430
rect 79382 400 79434 430
rect 79550 400 79602 430
rect 79718 400 79770 430
rect 79886 400 79938 430
rect 80054 400 80106 430
rect 80222 400 80274 430
rect 80390 400 80442 430
rect 80558 400 80610 430
rect 80726 400 80778 430
rect 80894 400 80946 430
rect 81062 400 81114 430
rect 81230 400 81282 430
rect 81398 400 81450 430
rect 81566 400 81618 430
rect 81734 400 81786 430
rect 81902 400 81954 430
rect 82070 400 82122 430
rect 82238 400 82290 430
rect 82406 400 82458 430
rect 82574 400 82626 430
rect 82742 400 82794 430
rect 82910 400 82962 430
rect 83078 400 83130 430
rect 83246 400 83298 430
rect 83414 400 83466 430
rect 83582 400 83634 430
rect 83750 400 83802 430
rect 83918 400 83970 430
rect 84086 400 84138 430
rect 84254 400 84306 430
rect 84422 400 84474 430
rect 84590 400 84642 430
rect 84758 400 84810 430
rect 84926 400 84978 430
rect 85094 400 85146 430
rect 85262 400 85314 430
rect 85430 400 85482 430
rect 85598 400 85650 430
rect 85766 400 85818 430
rect 85934 400 85986 430
rect 86102 400 86850 430
<< obsm3 >>
rect 2233 1554 86855 58898
<< metal4 >>
rect 2224 1538 2384 58438
rect 9904 1538 10064 58438
rect 17584 1538 17744 58438
rect 25264 1538 25424 58438
rect 32944 1538 33104 58438
rect 40624 1538 40784 58438
rect 48304 1538 48464 58438
rect 55984 1538 56144 58438
rect 63664 1538 63824 58438
rect 71344 1538 71504 58438
rect 79024 1538 79184 58438
rect 86704 1538 86864 58438
<< obsm4 >>
rect 53270 56793 55954 58063
rect 56174 56793 63042 58063
<< labels >>
rlabel metal2 s 3472 59600 3528 60000 6 io_active
port 1 nsew signal input
rlabel metal2 s 4200 59600 4256 60000 6 io_in[0]
port 2 nsew signal input
rlabel metal2 s 26040 59600 26096 60000 6 io_in[10]
port 3 nsew signal input
rlabel metal2 s 28224 59600 28280 60000 6 io_in[11]
port 4 nsew signal input
rlabel metal2 s 30408 59600 30464 60000 6 io_in[12]
port 5 nsew signal input
rlabel metal2 s 32592 59600 32648 60000 6 io_in[13]
port 6 nsew signal input
rlabel metal2 s 34776 59600 34832 60000 6 io_in[14]
port 7 nsew signal input
rlabel metal2 s 36960 59600 37016 60000 6 io_in[15]
port 8 nsew signal input
rlabel metal2 s 39144 59600 39200 60000 6 io_in[16]
port 9 nsew signal input
rlabel metal2 s 41328 59600 41384 60000 6 io_in[17]
port 10 nsew signal input
rlabel metal2 s 43512 59600 43568 60000 6 io_in[18]
port 11 nsew signal input
rlabel metal2 s 45696 59600 45752 60000 6 io_in[19]
port 12 nsew signal input
rlabel metal2 s 6384 59600 6440 60000 6 io_in[1]
port 13 nsew signal input
rlabel metal2 s 47880 59600 47936 60000 6 io_in[20]
port 14 nsew signal input
rlabel metal2 s 50064 59600 50120 60000 6 io_in[21]
port 15 nsew signal input
rlabel metal2 s 52248 59600 52304 60000 6 io_in[22]
port 16 nsew signal input
rlabel metal2 s 54432 59600 54488 60000 6 io_in[23]
port 17 nsew signal input
rlabel metal2 s 56616 59600 56672 60000 6 io_in[24]
port 18 nsew signal input
rlabel metal2 s 58800 59600 58856 60000 6 io_in[25]
port 19 nsew signal input
rlabel metal2 s 60984 59600 61040 60000 6 io_in[26]
port 20 nsew signal input
rlabel metal2 s 63168 59600 63224 60000 6 io_in[27]
port 21 nsew signal input
rlabel metal2 s 65352 59600 65408 60000 6 io_in[28]
port 22 nsew signal input
rlabel metal2 s 67536 59600 67592 60000 6 io_in[29]
port 23 nsew signal input
rlabel metal2 s 8568 59600 8624 60000 6 io_in[2]
port 24 nsew signal input
rlabel metal2 s 69720 59600 69776 60000 6 io_in[30]
port 25 nsew signal input
rlabel metal2 s 71904 59600 71960 60000 6 io_in[31]
port 26 nsew signal input
rlabel metal2 s 74088 59600 74144 60000 6 io_in[32]
port 27 nsew signal input
rlabel metal2 s 76272 59600 76328 60000 6 io_in[33]
port 28 nsew signal input
rlabel metal2 s 78456 59600 78512 60000 6 io_in[34]
port 29 nsew signal input
rlabel metal2 s 80640 59600 80696 60000 6 io_in[35]
port 30 nsew signal input
rlabel metal2 s 82824 59600 82880 60000 6 io_in[36]
port 31 nsew signal input
rlabel metal2 s 85008 59600 85064 60000 6 io_in[37]
port 32 nsew signal input
rlabel metal2 s 10752 59600 10808 60000 6 io_in[3]
port 33 nsew signal input
rlabel metal2 s 12936 59600 12992 60000 6 io_in[4]
port 34 nsew signal input
rlabel metal2 s 15120 59600 15176 60000 6 io_in[5]
port 35 nsew signal input
rlabel metal2 s 17304 59600 17360 60000 6 io_in[6]
port 36 nsew signal input
rlabel metal2 s 19488 59600 19544 60000 6 io_in[7]
port 37 nsew signal input
rlabel metal2 s 21672 59600 21728 60000 6 io_in[8]
port 38 nsew signal input
rlabel metal2 s 23856 59600 23912 60000 6 io_in[9]
port 39 nsew signal input
rlabel metal2 s 4928 59600 4984 60000 6 io_oeb[0]
port 40 nsew signal output
rlabel metal2 s 26768 59600 26824 60000 6 io_oeb[10]
port 41 nsew signal output
rlabel metal2 s 28952 59600 29008 60000 6 io_oeb[11]
port 42 nsew signal output
rlabel metal2 s 31136 59600 31192 60000 6 io_oeb[12]
port 43 nsew signal output
rlabel metal2 s 33320 59600 33376 60000 6 io_oeb[13]
port 44 nsew signal output
rlabel metal2 s 35504 59600 35560 60000 6 io_oeb[14]
port 45 nsew signal output
rlabel metal2 s 37688 59600 37744 60000 6 io_oeb[15]
port 46 nsew signal output
rlabel metal2 s 39872 59600 39928 60000 6 io_oeb[16]
port 47 nsew signal output
rlabel metal2 s 42056 59600 42112 60000 6 io_oeb[17]
port 48 nsew signal output
rlabel metal2 s 44240 59600 44296 60000 6 io_oeb[18]
port 49 nsew signal output
rlabel metal2 s 46424 59600 46480 60000 6 io_oeb[19]
port 50 nsew signal output
rlabel metal2 s 7112 59600 7168 60000 6 io_oeb[1]
port 51 nsew signal output
rlabel metal2 s 48608 59600 48664 60000 6 io_oeb[20]
port 52 nsew signal output
rlabel metal2 s 50792 59600 50848 60000 6 io_oeb[21]
port 53 nsew signal output
rlabel metal2 s 52976 59600 53032 60000 6 io_oeb[22]
port 54 nsew signal output
rlabel metal2 s 55160 59600 55216 60000 6 io_oeb[23]
port 55 nsew signal output
rlabel metal2 s 57344 59600 57400 60000 6 io_oeb[24]
port 56 nsew signal output
rlabel metal2 s 59528 59600 59584 60000 6 io_oeb[25]
port 57 nsew signal output
rlabel metal2 s 61712 59600 61768 60000 6 io_oeb[26]
port 58 nsew signal output
rlabel metal2 s 63896 59600 63952 60000 6 io_oeb[27]
port 59 nsew signal output
rlabel metal2 s 66080 59600 66136 60000 6 io_oeb[28]
port 60 nsew signal output
rlabel metal2 s 68264 59600 68320 60000 6 io_oeb[29]
port 61 nsew signal output
rlabel metal2 s 9296 59600 9352 60000 6 io_oeb[2]
port 62 nsew signal output
rlabel metal2 s 70448 59600 70504 60000 6 io_oeb[30]
port 63 nsew signal output
rlabel metal2 s 72632 59600 72688 60000 6 io_oeb[31]
port 64 nsew signal output
rlabel metal2 s 74816 59600 74872 60000 6 io_oeb[32]
port 65 nsew signal output
rlabel metal2 s 77000 59600 77056 60000 6 io_oeb[33]
port 66 nsew signal output
rlabel metal2 s 79184 59600 79240 60000 6 io_oeb[34]
port 67 nsew signal output
rlabel metal2 s 81368 59600 81424 60000 6 io_oeb[35]
port 68 nsew signal output
rlabel metal2 s 83552 59600 83608 60000 6 io_oeb[36]
port 69 nsew signal output
rlabel metal2 s 85736 59600 85792 60000 6 io_oeb[37]
port 70 nsew signal output
rlabel metal2 s 11480 59600 11536 60000 6 io_oeb[3]
port 71 nsew signal output
rlabel metal2 s 13664 59600 13720 60000 6 io_oeb[4]
port 72 nsew signal output
rlabel metal2 s 15848 59600 15904 60000 6 io_oeb[5]
port 73 nsew signal output
rlabel metal2 s 18032 59600 18088 60000 6 io_oeb[6]
port 74 nsew signal output
rlabel metal2 s 20216 59600 20272 60000 6 io_oeb[7]
port 75 nsew signal output
rlabel metal2 s 22400 59600 22456 60000 6 io_oeb[8]
port 76 nsew signal output
rlabel metal2 s 24584 59600 24640 60000 6 io_oeb[9]
port 77 nsew signal output
rlabel metal2 s 5656 59600 5712 60000 6 io_out[0]
port 78 nsew signal output
rlabel metal2 s 27496 59600 27552 60000 6 io_out[10]
port 79 nsew signal output
rlabel metal2 s 29680 59600 29736 60000 6 io_out[11]
port 80 nsew signal output
rlabel metal2 s 31864 59600 31920 60000 6 io_out[12]
port 81 nsew signal output
rlabel metal2 s 34048 59600 34104 60000 6 io_out[13]
port 82 nsew signal output
rlabel metal2 s 36232 59600 36288 60000 6 io_out[14]
port 83 nsew signal output
rlabel metal2 s 38416 59600 38472 60000 6 io_out[15]
port 84 nsew signal output
rlabel metal2 s 40600 59600 40656 60000 6 io_out[16]
port 85 nsew signal output
rlabel metal2 s 42784 59600 42840 60000 6 io_out[17]
port 86 nsew signal output
rlabel metal2 s 44968 59600 45024 60000 6 io_out[18]
port 87 nsew signal output
rlabel metal2 s 47152 59600 47208 60000 6 io_out[19]
port 88 nsew signal output
rlabel metal2 s 7840 59600 7896 60000 6 io_out[1]
port 89 nsew signal output
rlabel metal2 s 49336 59600 49392 60000 6 io_out[20]
port 90 nsew signal output
rlabel metal2 s 51520 59600 51576 60000 6 io_out[21]
port 91 nsew signal output
rlabel metal2 s 53704 59600 53760 60000 6 io_out[22]
port 92 nsew signal output
rlabel metal2 s 55888 59600 55944 60000 6 io_out[23]
port 93 nsew signal output
rlabel metal2 s 58072 59600 58128 60000 6 io_out[24]
port 94 nsew signal output
rlabel metal2 s 60256 59600 60312 60000 6 io_out[25]
port 95 nsew signal output
rlabel metal2 s 62440 59600 62496 60000 6 io_out[26]
port 96 nsew signal output
rlabel metal2 s 64624 59600 64680 60000 6 io_out[27]
port 97 nsew signal output
rlabel metal2 s 66808 59600 66864 60000 6 io_out[28]
port 98 nsew signal output
rlabel metal2 s 68992 59600 69048 60000 6 io_out[29]
port 99 nsew signal output
rlabel metal2 s 10024 59600 10080 60000 6 io_out[2]
port 100 nsew signal output
rlabel metal2 s 71176 59600 71232 60000 6 io_out[30]
port 101 nsew signal output
rlabel metal2 s 73360 59600 73416 60000 6 io_out[31]
port 102 nsew signal output
rlabel metal2 s 75544 59600 75600 60000 6 io_out[32]
port 103 nsew signal output
rlabel metal2 s 77728 59600 77784 60000 6 io_out[33]
port 104 nsew signal output
rlabel metal2 s 79912 59600 79968 60000 6 io_out[34]
port 105 nsew signal output
rlabel metal2 s 82096 59600 82152 60000 6 io_out[35]
port 106 nsew signal output
rlabel metal2 s 84280 59600 84336 60000 6 io_out[36]
port 107 nsew signal output
rlabel metal2 s 86464 59600 86520 60000 6 io_out[37]
port 108 nsew signal output
rlabel metal2 s 12208 59600 12264 60000 6 io_out[3]
port 109 nsew signal output
rlabel metal2 s 14392 59600 14448 60000 6 io_out[4]
port 110 nsew signal output
rlabel metal2 s 16576 59600 16632 60000 6 io_out[5]
port 111 nsew signal output
rlabel metal2 s 18760 59600 18816 60000 6 io_out[6]
port 112 nsew signal output
rlabel metal2 s 20944 59600 21000 60000 6 io_out[7]
port 113 nsew signal output
rlabel metal2 s 23128 59600 23184 60000 6 io_out[8]
port 114 nsew signal output
rlabel metal2 s 25312 59600 25368 60000 6 io_out[9]
port 115 nsew signal output
rlabel metal2 s 21672 0 21728 400 6 la_data_in[0]
port 116 nsew signal input
rlabel metal2 s 72072 0 72128 400 6 la_data_in[100]
port 117 nsew signal input
rlabel metal2 s 72576 0 72632 400 6 la_data_in[101]
port 118 nsew signal input
rlabel metal2 s 73080 0 73136 400 6 la_data_in[102]
port 119 nsew signal input
rlabel metal2 s 73584 0 73640 400 6 la_data_in[103]
port 120 nsew signal input
rlabel metal2 s 74088 0 74144 400 6 la_data_in[104]
port 121 nsew signal input
rlabel metal2 s 74592 0 74648 400 6 la_data_in[105]
port 122 nsew signal input
rlabel metal2 s 75096 0 75152 400 6 la_data_in[106]
port 123 nsew signal input
rlabel metal2 s 75600 0 75656 400 6 la_data_in[107]
port 124 nsew signal input
rlabel metal2 s 76104 0 76160 400 6 la_data_in[108]
port 125 nsew signal input
rlabel metal2 s 76608 0 76664 400 6 la_data_in[109]
port 126 nsew signal input
rlabel metal2 s 26712 0 26768 400 6 la_data_in[10]
port 127 nsew signal input
rlabel metal2 s 77112 0 77168 400 6 la_data_in[110]
port 128 nsew signal input
rlabel metal2 s 77616 0 77672 400 6 la_data_in[111]
port 129 nsew signal input
rlabel metal2 s 78120 0 78176 400 6 la_data_in[112]
port 130 nsew signal input
rlabel metal2 s 78624 0 78680 400 6 la_data_in[113]
port 131 nsew signal input
rlabel metal2 s 79128 0 79184 400 6 la_data_in[114]
port 132 nsew signal input
rlabel metal2 s 79632 0 79688 400 6 la_data_in[115]
port 133 nsew signal input
rlabel metal2 s 80136 0 80192 400 6 la_data_in[116]
port 134 nsew signal input
rlabel metal2 s 80640 0 80696 400 6 la_data_in[117]
port 135 nsew signal input
rlabel metal2 s 81144 0 81200 400 6 la_data_in[118]
port 136 nsew signal input
rlabel metal2 s 81648 0 81704 400 6 la_data_in[119]
port 137 nsew signal input
rlabel metal2 s 27216 0 27272 400 6 la_data_in[11]
port 138 nsew signal input
rlabel metal2 s 82152 0 82208 400 6 la_data_in[120]
port 139 nsew signal input
rlabel metal2 s 82656 0 82712 400 6 la_data_in[121]
port 140 nsew signal input
rlabel metal2 s 83160 0 83216 400 6 la_data_in[122]
port 141 nsew signal input
rlabel metal2 s 83664 0 83720 400 6 la_data_in[123]
port 142 nsew signal input
rlabel metal2 s 84168 0 84224 400 6 la_data_in[124]
port 143 nsew signal input
rlabel metal2 s 84672 0 84728 400 6 la_data_in[125]
port 144 nsew signal input
rlabel metal2 s 85176 0 85232 400 6 la_data_in[126]
port 145 nsew signal input
rlabel metal2 s 85680 0 85736 400 6 la_data_in[127]
port 146 nsew signal input
rlabel metal2 s 27720 0 27776 400 6 la_data_in[12]
port 147 nsew signal input
rlabel metal2 s 28224 0 28280 400 6 la_data_in[13]
port 148 nsew signal input
rlabel metal2 s 28728 0 28784 400 6 la_data_in[14]
port 149 nsew signal input
rlabel metal2 s 29232 0 29288 400 6 la_data_in[15]
port 150 nsew signal input
rlabel metal2 s 29736 0 29792 400 6 la_data_in[16]
port 151 nsew signal input
rlabel metal2 s 30240 0 30296 400 6 la_data_in[17]
port 152 nsew signal input
rlabel metal2 s 30744 0 30800 400 6 la_data_in[18]
port 153 nsew signal input
rlabel metal2 s 31248 0 31304 400 6 la_data_in[19]
port 154 nsew signal input
rlabel metal2 s 22176 0 22232 400 6 la_data_in[1]
port 155 nsew signal input
rlabel metal2 s 31752 0 31808 400 6 la_data_in[20]
port 156 nsew signal input
rlabel metal2 s 32256 0 32312 400 6 la_data_in[21]
port 157 nsew signal input
rlabel metal2 s 32760 0 32816 400 6 la_data_in[22]
port 158 nsew signal input
rlabel metal2 s 33264 0 33320 400 6 la_data_in[23]
port 159 nsew signal input
rlabel metal2 s 33768 0 33824 400 6 la_data_in[24]
port 160 nsew signal input
rlabel metal2 s 34272 0 34328 400 6 la_data_in[25]
port 161 nsew signal input
rlabel metal2 s 34776 0 34832 400 6 la_data_in[26]
port 162 nsew signal input
rlabel metal2 s 35280 0 35336 400 6 la_data_in[27]
port 163 nsew signal input
rlabel metal2 s 35784 0 35840 400 6 la_data_in[28]
port 164 nsew signal input
rlabel metal2 s 36288 0 36344 400 6 la_data_in[29]
port 165 nsew signal input
rlabel metal2 s 22680 0 22736 400 6 la_data_in[2]
port 166 nsew signal input
rlabel metal2 s 36792 0 36848 400 6 la_data_in[30]
port 167 nsew signal input
rlabel metal2 s 37296 0 37352 400 6 la_data_in[31]
port 168 nsew signal input
rlabel metal2 s 37800 0 37856 400 6 la_data_in[32]
port 169 nsew signal input
rlabel metal2 s 38304 0 38360 400 6 la_data_in[33]
port 170 nsew signal input
rlabel metal2 s 38808 0 38864 400 6 la_data_in[34]
port 171 nsew signal input
rlabel metal2 s 39312 0 39368 400 6 la_data_in[35]
port 172 nsew signal input
rlabel metal2 s 39816 0 39872 400 6 la_data_in[36]
port 173 nsew signal input
rlabel metal2 s 40320 0 40376 400 6 la_data_in[37]
port 174 nsew signal input
rlabel metal2 s 40824 0 40880 400 6 la_data_in[38]
port 175 nsew signal input
rlabel metal2 s 41328 0 41384 400 6 la_data_in[39]
port 176 nsew signal input
rlabel metal2 s 23184 0 23240 400 6 la_data_in[3]
port 177 nsew signal input
rlabel metal2 s 41832 0 41888 400 6 la_data_in[40]
port 178 nsew signal input
rlabel metal2 s 42336 0 42392 400 6 la_data_in[41]
port 179 nsew signal input
rlabel metal2 s 42840 0 42896 400 6 la_data_in[42]
port 180 nsew signal input
rlabel metal2 s 43344 0 43400 400 6 la_data_in[43]
port 181 nsew signal input
rlabel metal2 s 43848 0 43904 400 6 la_data_in[44]
port 182 nsew signal input
rlabel metal2 s 44352 0 44408 400 6 la_data_in[45]
port 183 nsew signal input
rlabel metal2 s 44856 0 44912 400 6 la_data_in[46]
port 184 nsew signal input
rlabel metal2 s 45360 0 45416 400 6 la_data_in[47]
port 185 nsew signal input
rlabel metal2 s 45864 0 45920 400 6 la_data_in[48]
port 186 nsew signal input
rlabel metal2 s 46368 0 46424 400 6 la_data_in[49]
port 187 nsew signal input
rlabel metal2 s 23688 0 23744 400 6 la_data_in[4]
port 188 nsew signal input
rlabel metal2 s 46872 0 46928 400 6 la_data_in[50]
port 189 nsew signal input
rlabel metal2 s 47376 0 47432 400 6 la_data_in[51]
port 190 nsew signal input
rlabel metal2 s 47880 0 47936 400 6 la_data_in[52]
port 191 nsew signal input
rlabel metal2 s 48384 0 48440 400 6 la_data_in[53]
port 192 nsew signal input
rlabel metal2 s 48888 0 48944 400 6 la_data_in[54]
port 193 nsew signal input
rlabel metal2 s 49392 0 49448 400 6 la_data_in[55]
port 194 nsew signal input
rlabel metal2 s 49896 0 49952 400 6 la_data_in[56]
port 195 nsew signal input
rlabel metal2 s 50400 0 50456 400 6 la_data_in[57]
port 196 nsew signal input
rlabel metal2 s 50904 0 50960 400 6 la_data_in[58]
port 197 nsew signal input
rlabel metal2 s 51408 0 51464 400 6 la_data_in[59]
port 198 nsew signal input
rlabel metal2 s 24192 0 24248 400 6 la_data_in[5]
port 199 nsew signal input
rlabel metal2 s 51912 0 51968 400 6 la_data_in[60]
port 200 nsew signal input
rlabel metal2 s 52416 0 52472 400 6 la_data_in[61]
port 201 nsew signal input
rlabel metal2 s 52920 0 52976 400 6 la_data_in[62]
port 202 nsew signal input
rlabel metal2 s 53424 0 53480 400 6 la_data_in[63]
port 203 nsew signal input
rlabel metal2 s 53928 0 53984 400 6 la_data_in[64]
port 204 nsew signal input
rlabel metal2 s 54432 0 54488 400 6 la_data_in[65]
port 205 nsew signal input
rlabel metal2 s 54936 0 54992 400 6 la_data_in[66]
port 206 nsew signal input
rlabel metal2 s 55440 0 55496 400 6 la_data_in[67]
port 207 nsew signal input
rlabel metal2 s 55944 0 56000 400 6 la_data_in[68]
port 208 nsew signal input
rlabel metal2 s 56448 0 56504 400 6 la_data_in[69]
port 209 nsew signal input
rlabel metal2 s 24696 0 24752 400 6 la_data_in[6]
port 210 nsew signal input
rlabel metal2 s 56952 0 57008 400 6 la_data_in[70]
port 211 nsew signal input
rlabel metal2 s 57456 0 57512 400 6 la_data_in[71]
port 212 nsew signal input
rlabel metal2 s 57960 0 58016 400 6 la_data_in[72]
port 213 nsew signal input
rlabel metal2 s 58464 0 58520 400 6 la_data_in[73]
port 214 nsew signal input
rlabel metal2 s 58968 0 59024 400 6 la_data_in[74]
port 215 nsew signal input
rlabel metal2 s 59472 0 59528 400 6 la_data_in[75]
port 216 nsew signal input
rlabel metal2 s 59976 0 60032 400 6 la_data_in[76]
port 217 nsew signal input
rlabel metal2 s 60480 0 60536 400 6 la_data_in[77]
port 218 nsew signal input
rlabel metal2 s 60984 0 61040 400 6 la_data_in[78]
port 219 nsew signal input
rlabel metal2 s 61488 0 61544 400 6 la_data_in[79]
port 220 nsew signal input
rlabel metal2 s 25200 0 25256 400 6 la_data_in[7]
port 221 nsew signal input
rlabel metal2 s 61992 0 62048 400 6 la_data_in[80]
port 222 nsew signal input
rlabel metal2 s 62496 0 62552 400 6 la_data_in[81]
port 223 nsew signal input
rlabel metal2 s 63000 0 63056 400 6 la_data_in[82]
port 224 nsew signal input
rlabel metal2 s 63504 0 63560 400 6 la_data_in[83]
port 225 nsew signal input
rlabel metal2 s 64008 0 64064 400 6 la_data_in[84]
port 226 nsew signal input
rlabel metal2 s 64512 0 64568 400 6 la_data_in[85]
port 227 nsew signal input
rlabel metal2 s 65016 0 65072 400 6 la_data_in[86]
port 228 nsew signal input
rlabel metal2 s 65520 0 65576 400 6 la_data_in[87]
port 229 nsew signal input
rlabel metal2 s 66024 0 66080 400 6 la_data_in[88]
port 230 nsew signal input
rlabel metal2 s 66528 0 66584 400 6 la_data_in[89]
port 231 nsew signal input
rlabel metal2 s 25704 0 25760 400 6 la_data_in[8]
port 232 nsew signal input
rlabel metal2 s 67032 0 67088 400 6 la_data_in[90]
port 233 nsew signal input
rlabel metal2 s 67536 0 67592 400 6 la_data_in[91]
port 234 nsew signal input
rlabel metal2 s 68040 0 68096 400 6 la_data_in[92]
port 235 nsew signal input
rlabel metal2 s 68544 0 68600 400 6 la_data_in[93]
port 236 nsew signal input
rlabel metal2 s 69048 0 69104 400 6 la_data_in[94]
port 237 nsew signal input
rlabel metal2 s 69552 0 69608 400 6 la_data_in[95]
port 238 nsew signal input
rlabel metal2 s 70056 0 70112 400 6 la_data_in[96]
port 239 nsew signal input
rlabel metal2 s 70560 0 70616 400 6 la_data_in[97]
port 240 nsew signal input
rlabel metal2 s 71064 0 71120 400 6 la_data_in[98]
port 241 nsew signal input
rlabel metal2 s 71568 0 71624 400 6 la_data_in[99]
port 242 nsew signal input
rlabel metal2 s 26208 0 26264 400 6 la_data_in[9]
port 243 nsew signal input
rlabel metal2 s 21840 0 21896 400 6 la_data_out[0]
port 244 nsew signal output
rlabel metal2 s 72240 0 72296 400 6 la_data_out[100]
port 245 nsew signal output
rlabel metal2 s 72744 0 72800 400 6 la_data_out[101]
port 246 nsew signal output
rlabel metal2 s 73248 0 73304 400 6 la_data_out[102]
port 247 nsew signal output
rlabel metal2 s 73752 0 73808 400 6 la_data_out[103]
port 248 nsew signal output
rlabel metal2 s 74256 0 74312 400 6 la_data_out[104]
port 249 nsew signal output
rlabel metal2 s 74760 0 74816 400 6 la_data_out[105]
port 250 nsew signal output
rlabel metal2 s 75264 0 75320 400 6 la_data_out[106]
port 251 nsew signal output
rlabel metal2 s 75768 0 75824 400 6 la_data_out[107]
port 252 nsew signal output
rlabel metal2 s 76272 0 76328 400 6 la_data_out[108]
port 253 nsew signal output
rlabel metal2 s 76776 0 76832 400 6 la_data_out[109]
port 254 nsew signal output
rlabel metal2 s 26880 0 26936 400 6 la_data_out[10]
port 255 nsew signal output
rlabel metal2 s 77280 0 77336 400 6 la_data_out[110]
port 256 nsew signal output
rlabel metal2 s 77784 0 77840 400 6 la_data_out[111]
port 257 nsew signal output
rlabel metal2 s 78288 0 78344 400 6 la_data_out[112]
port 258 nsew signal output
rlabel metal2 s 78792 0 78848 400 6 la_data_out[113]
port 259 nsew signal output
rlabel metal2 s 79296 0 79352 400 6 la_data_out[114]
port 260 nsew signal output
rlabel metal2 s 79800 0 79856 400 6 la_data_out[115]
port 261 nsew signal output
rlabel metal2 s 80304 0 80360 400 6 la_data_out[116]
port 262 nsew signal output
rlabel metal2 s 80808 0 80864 400 6 la_data_out[117]
port 263 nsew signal output
rlabel metal2 s 81312 0 81368 400 6 la_data_out[118]
port 264 nsew signal output
rlabel metal2 s 81816 0 81872 400 6 la_data_out[119]
port 265 nsew signal output
rlabel metal2 s 27384 0 27440 400 6 la_data_out[11]
port 266 nsew signal output
rlabel metal2 s 82320 0 82376 400 6 la_data_out[120]
port 267 nsew signal output
rlabel metal2 s 82824 0 82880 400 6 la_data_out[121]
port 268 nsew signal output
rlabel metal2 s 83328 0 83384 400 6 la_data_out[122]
port 269 nsew signal output
rlabel metal2 s 83832 0 83888 400 6 la_data_out[123]
port 270 nsew signal output
rlabel metal2 s 84336 0 84392 400 6 la_data_out[124]
port 271 nsew signal output
rlabel metal2 s 84840 0 84896 400 6 la_data_out[125]
port 272 nsew signal output
rlabel metal2 s 85344 0 85400 400 6 la_data_out[126]
port 273 nsew signal output
rlabel metal2 s 85848 0 85904 400 6 la_data_out[127]
port 274 nsew signal output
rlabel metal2 s 27888 0 27944 400 6 la_data_out[12]
port 275 nsew signal output
rlabel metal2 s 28392 0 28448 400 6 la_data_out[13]
port 276 nsew signal output
rlabel metal2 s 28896 0 28952 400 6 la_data_out[14]
port 277 nsew signal output
rlabel metal2 s 29400 0 29456 400 6 la_data_out[15]
port 278 nsew signal output
rlabel metal2 s 29904 0 29960 400 6 la_data_out[16]
port 279 nsew signal output
rlabel metal2 s 30408 0 30464 400 6 la_data_out[17]
port 280 nsew signal output
rlabel metal2 s 30912 0 30968 400 6 la_data_out[18]
port 281 nsew signal output
rlabel metal2 s 31416 0 31472 400 6 la_data_out[19]
port 282 nsew signal output
rlabel metal2 s 22344 0 22400 400 6 la_data_out[1]
port 283 nsew signal output
rlabel metal2 s 31920 0 31976 400 6 la_data_out[20]
port 284 nsew signal output
rlabel metal2 s 32424 0 32480 400 6 la_data_out[21]
port 285 nsew signal output
rlabel metal2 s 32928 0 32984 400 6 la_data_out[22]
port 286 nsew signal output
rlabel metal2 s 33432 0 33488 400 6 la_data_out[23]
port 287 nsew signal output
rlabel metal2 s 33936 0 33992 400 6 la_data_out[24]
port 288 nsew signal output
rlabel metal2 s 34440 0 34496 400 6 la_data_out[25]
port 289 nsew signal output
rlabel metal2 s 34944 0 35000 400 6 la_data_out[26]
port 290 nsew signal output
rlabel metal2 s 35448 0 35504 400 6 la_data_out[27]
port 291 nsew signal output
rlabel metal2 s 35952 0 36008 400 6 la_data_out[28]
port 292 nsew signal output
rlabel metal2 s 36456 0 36512 400 6 la_data_out[29]
port 293 nsew signal output
rlabel metal2 s 22848 0 22904 400 6 la_data_out[2]
port 294 nsew signal output
rlabel metal2 s 36960 0 37016 400 6 la_data_out[30]
port 295 nsew signal output
rlabel metal2 s 37464 0 37520 400 6 la_data_out[31]
port 296 nsew signal output
rlabel metal2 s 37968 0 38024 400 6 la_data_out[32]
port 297 nsew signal output
rlabel metal2 s 38472 0 38528 400 6 la_data_out[33]
port 298 nsew signal output
rlabel metal2 s 38976 0 39032 400 6 la_data_out[34]
port 299 nsew signal output
rlabel metal2 s 39480 0 39536 400 6 la_data_out[35]
port 300 nsew signal output
rlabel metal2 s 39984 0 40040 400 6 la_data_out[36]
port 301 nsew signal output
rlabel metal2 s 40488 0 40544 400 6 la_data_out[37]
port 302 nsew signal output
rlabel metal2 s 40992 0 41048 400 6 la_data_out[38]
port 303 nsew signal output
rlabel metal2 s 41496 0 41552 400 6 la_data_out[39]
port 304 nsew signal output
rlabel metal2 s 23352 0 23408 400 6 la_data_out[3]
port 305 nsew signal output
rlabel metal2 s 42000 0 42056 400 6 la_data_out[40]
port 306 nsew signal output
rlabel metal2 s 42504 0 42560 400 6 la_data_out[41]
port 307 nsew signal output
rlabel metal2 s 43008 0 43064 400 6 la_data_out[42]
port 308 nsew signal output
rlabel metal2 s 43512 0 43568 400 6 la_data_out[43]
port 309 nsew signal output
rlabel metal2 s 44016 0 44072 400 6 la_data_out[44]
port 310 nsew signal output
rlabel metal2 s 44520 0 44576 400 6 la_data_out[45]
port 311 nsew signal output
rlabel metal2 s 45024 0 45080 400 6 la_data_out[46]
port 312 nsew signal output
rlabel metal2 s 45528 0 45584 400 6 la_data_out[47]
port 313 nsew signal output
rlabel metal2 s 46032 0 46088 400 6 la_data_out[48]
port 314 nsew signal output
rlabel metal2 s 46536 0 46592 400 6 la_data_out[49]
port 315 nsew signal output
rlabel metal2 s 23856 0 23912 400 6 la_data_out[4]
port 316 nsew signal output
rlabel metal2 s 47040 0 47096 400 6 la_data_out[50]
port 317 nsew signal output
rlabel metal2 s 47544 0 47600 400 6 la_data_out[51]
port 318 nsew signal output
rlabel metal2 s 48048 0 48104 400 6 la_data_out[52]
port 319 nsew signal output
rlabel metal2 s 48552 0 48608 400 6 la_data_out[53]
port 320 nsew signal output
rlabel metal2 s 49056 0 49112 400 6 la_data_out[54]
port 321 nsew signal output
rlabel metal2 s 49560 0 49616 400 6 la_data_out[55]
port 322 nsew signal output
rlabel metal2 s 50064 0 50120 400 6 la_data_out[56]
port 323 nsew signal output
rlabel metal2 s 50568 0 50624 400 6 la_data_out[57]
port 324 nsew signal output
rlabel metal2 s 51072 0 51128 400 6 la_data_out[58]
port 325 nsew signal output
rlabel metal2 s 51576 0 51632 400 6 la_data_out[59]
port 326 nsew signal output
rlabel metal2 s 24360 0 24416 400 6 la_data_out[5]
port 327 nsew signal output
rlabel metal2 s 52080 0 52136 400 6 la_data_out[60]
port 328 nsew signal output
rlabel metal2 s 52584 0 52640 400 6 la_data_out[61]
port 329 nsew signal output
rlabel metal2 s 53088 0 53144 400 6 la_data_out[62]
port 330 nsew signal output
rlabel metal2 s 53592 0 53648 400 6 la_data_out[63]
port 331 nsew signal output
rlabel metal2 s 54096 0 54152 400 6 la_data_out[64]
port 332 nsew signal output
rlabel metal2 s 54600 0 54656 400 6 la_data_out[65]
port 333 nsew signal output
rlabel metal2 s 55104 0 55160 400 6 la_data_out[66]
port 334 nsew signal output
rlabel metal2 s 55608 0 55664 400 6 la_data_out[67]
port 335 nsew signal output
rlabel metal2 s 56112 0 56168 400 6 la_data_out[68]
port 336 nsew signal output
rlabel metal2 s 56616 0 56672 400 6 la_data_out[69]
port 337 nsew signal output
rlabel metal2 s 24864 0 24920 400 6 la_data_out[6]
port 338 nsew signal output
rlabel metal2 s 57120 0 57176 400 6 la_data_out[70]
port 339 nsew signal output
rlabel metal2 s 57624 0 57680 400 6 la_data_out[71]
port 340 nsew signal output
rlabel metal2 s 58128 0 58184 400 6 la_data_out[72]
port 341 nsew signal output
rlabel metal2 s 58632 0 58688 400 6 la_data_out[73]
port 342 nsew signal output
rlabel metal2 s 59136 0 59192 400 6 la_data_out[74]
port 343 nsew signal output
rlabel metal2 s 59640 0 59696 400 6 la_data_out[75]
port 344 nsew signal output
rlabel metal2 s 60144 0 60200 400 6 la_data_out[76]
port 345 nsew signal output
rlabel metal2 s 60648 0 60704 400 6 la_data_out[77]
port 346 nsew signal output
rlabel metal2 s 61152 0 61208 400 6 la_data_out[78]
port 347 nsew signal output
rlabel metal2 s 61656 0 61712 400 6 la_data_out[79]
port 348 nsew signal output
rlabel metal2 s 25368 0 25424 400 6 la_data_out[7]
port 349 nsew signal output
rlabel metal2 s 62160 0 62216 400 6 la_data_out[80]
port 350 nsew signal output
rlabel metal2 s 62664 0 62720 400 6 la_data_out[81]
port 351 nsew signal output
rlabel metal2 s 63168 0 63224 400 6 la_data_out[82]
port 352 nsew signal output
rlabel metal2 s 63672 0 63728 400 6 la_data_out[83]
port 353 nsew signal output
rlabel metal2 s 64176 0 64232 400 6 la_data_out[84]
port 354 nsew signal output
rlabel metal2 s 64680 0 64736 400 6 la_data_out[85]
port 355 nsew signal output
rlabel metal2 s 65184 0 65240 400 6 la_data_out[86]
port 356 nsew signal output
rlabel metal2 s 65688 0 65744 400 6 la_data_out[87]
port 357 nsew signal output
rlabel metal2 s 66192 0 66248 400 6 la_data_out[88]
port 358 nsew signal output
rlabel metal2 s 66696 0 66752 400 6 la_data_out[89]
port 359 nsew signal output
rlabel metal2 s 25872 0 25928 400 6 la_data_out[8]
port 360 nsew signal output
rlabel metal2 s 67200 0 67256 400 6 la_data_out[90]
port 361 nsew signal output
rlabel metal2 s 67704 0 67760 400 6 la_data_out[91]
port 362 nsew signal output
rlabel metal2 s 68208 0 68264 400 6 la_data_out[92]
port 363 nsew signal output
rlabel metal2 s 68712 0 68768 400 6 la_data_out[93]
port 364 nsew signal output
rlabel metal2 s 69216 0 69272 400 6 la_data_out[94]
port 365 nsew signal output
rlabel metal2 s 69720 0 69776 400 6 la_data_out[95]
port 366 nsew signal output
rlabel metal2 s 70224 0 70280 400 6 la_data_out[96]
port 367 nsew signal output
rlabel metal2 s 70728 0 70784 400 6 la_data_out[97]
port 368 nsew signal output
rlabel metal2 s 71232 0 71288 400 6 la_data_out[98]
port 369 nsew signal output
rlabel metal2 s 71736 0 71792 400 6 la_data_out[99]
port 370 nsew signal output
rlabel metal2 s 26376 0 26432 400 6 la_data_out[9]
port 371 nsew signal output
rlabel metal2 s 22008 0 22064 400 6 la_oenb[0]
port 372 nsew signal input
rlabel metal2 s 72408 0 72464 400 6 la_oenb[100]
port 373 nsew signal input
rlabel metal2 s 72912 0 72968 400 6 la_oenb[101]
port 374 nsew signal input
rlabel metal2 s 73416 0 73472 400 6 la_oenb[102]
port 375 nsew signal input
rlabel metal2 s 73920 0 73976 400 6 la_oenb[103]
port 376 nsew signal input
rlabel metal2 s 74424 0 74480 400 6 la_oenb[104]
port 377 nsew signal input
rlabel metal2 s 74928 0 74984 400 6 la_oenb[105]
port 378 nsew signal input
rlabel metal2 s 75432 0 75488 400 6 la_oenb[106]
port 379 nsew signal input
rlabel metal2 s 75936 0 75992 400 6 la_oenb[107]
port 380 nsew signal input
rlabel metal2 s 76440 0 76496 400 6 la_oenb[108]
port 381 nsew signal input
rlabel metal2 s 76944 0 77000 400 6 la_oenb[109]
port 382 nsew signal input
rlabel metal2 s 27048 0 27104 400 6 la_oenb[10]
port 383 nsew signal input
rlabel metal2 s 77448 0 77504 400 6 la_oenb[110]
port 384 nsew signal input
rlabel metal2 s 77952 0 78008 400 6 la_oenb[111]
port 385 nsew signal input
rlabel metal2 s 78456 0 78512 400 6 la_oenb[112]
port 386 nsew signal input
rlabel metal2 s 78960 0 79016 400 6 la_oenb[113]
port 387 nsew signal input
rlabel metal2 s 79464 0 79520 400 6 la_oenb[114]
port 388 nsew signal input
rlabel metal2 s 79968 0 80024 400 6 la_oenb[115]
port 389 nsew signal input
rlabel metal2 s 80472 0 80528 400 6 la_oenb[116]
port 390 nsew signal input
rlabel metal2 s 80976 0 81032 400 6 la_oenb[117]
port 391 nsew signal input
rlabel metal2 s 81480 0 81536 400 6 la_oenb[118]
port 392 nsew signal input
rlabel metal2 s 81984 0 82040 400 6 la_oenb[119]
port 393 nsew signal input
rlabel metal2 s 27552 0 27608 400 6 la_oenb[11]
port 394 nsew signal input
rlabel metal2 s 82488 0 82544 400 6 la_oenb[120]
port 395 nsew signal input
rlabel metal2 s 82992 0 83048 400 6 la_oenb[121]
port 396 nsew signal input
rlabel metal2 s 83496 0 83552 400 6 la_oenb[122]
port 397 nsew signal input
rlabel metal2 s 84000 0 84056 400 6 la_oenb[123]
port 398 nsew signal input
rlabel metal2 s 84504 0 84560 400 6 la_oenb[124]
port 399 nsew signal input
rlabel metal2 s 85008 0 85064 400 6 la_oenb[125]
port 400 nsew signal input
rlabel metal2 s 85512 0 85568 400 6 la_oenb[126]
port 401 nsew signal input
rlabel metal2 s 86016 0 86072 400 6 la_oenb[127]
port 402 nsew signal input
rlabel metal2 s 28056 0 28112 400 6 la_oenb[12]
port 403 nsew signal input
rlabel metal2 s 28560 0 28616 400 6 la_oenb[13]
port 404 nsew signal input
rlabel metal2 s 29064 0 29120 400 6 la_oenb[14]
port 405 nsew signal input
rlabel metal2 s 29568 0 29624 400 6 la_oenb[15]
port 406 nsew signal input
rlabel metal2 s 30072 0 30128 400 6 la_oenb[16]
port 407 nsew signal input
rlabel metal2 s 30576 0 30632 400 6 la_oenb[17]
port 408 nsew signal input
rlabel metal2 s 31080 0 31136 400 6 la_oenb[18]
port 409 nsew signal input
rlabel metal2 s 31584 0 31640 400 6 la_oenb[19]
port 410 nsew signal input
rlabel metal2 s 22512 0 22568 400 6 la_oenb[1]
port 411 nsew signal input
rlabel metal2 s 32088 0 32144 400 6 la_oenb[20]
port 412 nsew signal input
rlabel metal2 s 32592 0 32648 400 6 la_oenb[21]
port 413 nsew signal input
rlabel metal2 s 33096 0 33152 400 6 la_oenb[22]
port 414 nsew signal input
rlabel metal2 s 33600 0 33656 400 6 la_oenb[23]
port 415 nsew signal input
rlabel metal2 s 34104 0 34160 400 6 la_oenb[24]
port 416 nsew signal input
rlabel metal2 s 34608 0 34664 400 6 la_oenb[25]
port 417 nsew signal input
rlabel metal2 s 35112 0 35168 400 6 la_oenb[26]
port 418 nsew signal input
rlabel metal2 s 35616 0 35672 400 6 la_oenb[27]
port 419 nsew signal input
rlabel metal2 s 36120 0 36176 400 6 la_oenb[28]
port 420 nsew signal input
rlabel metal2 s 36624 0 36680 400 6 la_oenb[29]
port 421 nsew signal input
rlabel metal2 s 23016 0 23072 400 6 la_oenb[2]
port 422 nsew signal input
rlabel metal2 s 37128 0 37184 400 6 la_oenb[30]
port 423 nsew signal input
rlabel metal2 s 37632 0 37688 400 6 la_oenb[31]
port 424 nsew signal input
rlabel metal2 s 38136 0 38192 400 6 la_oenb[32]
port 425 nsew signal input
rlabel metal2 s 38640 0 38696 400 6 la_oenb[33]
port 426 nsew signal input
rlabel metal2 s 39144 0 39200 400 6 la_oenb[34]
port 427 nsew signal input
rlabel metal2 s 39648 0 39704 400 6 la_oenb[35]
port 428 nsew signal input
rlabel metal2 s 40152 0 40208 400 6 la_oenb[36]
port 429 nsew signal input
rlabel metal2 s 40656 0 40712 400 6 la_oenb[37]
port 430 nsew signal input
rlabel metal2 s 41160 0 41216 400 6 la_oenb[38]
port 431 nsew signal input
rlabel metal2 s 41664 0 41720 400 6 la_oenb[39]
port 432 nsew signal input
rlabel metal2 s 23520 0 23576 400 6 la_oenb[3]
port 433 nsew signal input
rlabel metal2 s 42168 0 42224 400 6 la_oenb[40]
port 434 nsew signal input
rlabel metal2 s 42672 0 42728 400 6 la_oenb[41]
port 435 nsew signal input
rlabel metal2 s 43176 0 43232 400 6 la_oenb[42]
port 436 nsew signal input
rlabel metal2 s 43680 0 43736 400 6 la_oenb[43]
port 437 nsew signal input
rlabel metal2 s 44184 0 44240 400 6 la_oenb[44]
port 438 nsew signal input
rlabel metal2 s 44688 0 44744 400 6 la_oenb[45]
port 439 nsew signal input
rlabel metal2 s 45192 0 45248 400 6 la_oenb[46]
port 440 nsew signal input
rlabel metal2 s 45696 0 45752 400 6 la_oenb[47]
port 441 nsew signal input
rlabel metal2 s 46200 0 46256 400 6 la_oenb[48]
port 442 nsew signal input
rlabel metal2 s 46704 0 46760 400 6 la_oenb[49]
port 443 nsew signal input
rlabel metal2 s 24024 0 24080 400 6 la_oenb[4]
port 444 nsew signal input
rlabel metal2 s 47208 0 47264 400 6 la_oenb[50]
port 445 nsew signal input
rlabel metal2 s 47712 0 47768 400 6 la_oenb[51]
port 446 nsew signal input
rlabel metal2 s 48216 0 48272 400 6 la_oenb[52]
port 447 nsew signal input
rlabel metal2 s 48720 0 48776 400 6 la_oenb[53]
port 448 nsew signal input
rlabel metal2 s 49224 0 49280 400 6 la_oenb[54]
port 449 nsew signal input
rlabel metal2 s 49728 0 49784 400 6 la_oenb[55]
port 450 nsew signal input
rlabel metal2 s 50232 0 50288 400 6 la_oenb[56]
port 451 nsew signal input
rlabel metal2 s 50736 0 50792 400 6 la_oenb[57]
port 452 nsew signal input
rlabel metal2 s 51240 0 51296 400 6 la_oenb[58]
port 453 nsew signal input
rlabel metal2 s 51744 0 51800 400 6 la_oenb[59]
port 454 nsew signal input
rlabel metal2 s 24528 0 24584 400 6 la_oenb[5]
port 455 nsew signal input
rlabel metal2 s 52248 0 52304 400 6 la_oenb[60]
port 456 nsew signal input
rlabel metal2 s 52752 0 52808 400 6 la_oenb[61]
port 457 nsew signal input
rlabel metal2 s 53256 0 53312 400 6 la_oenb[62]
port 458 nsew signal input
rlabel metal2 s 53760 0 53816 400 6 la_oenb[63]
port 459 nsew signal input
rlabel metal2 s 54264 0 54320 400 6 la_oenb[64]
port 460 nsew signal input
rlabel metal2 s 54768 0 54824 400 6 la_oenb[65]
port 461 nsew signal input
rlabel metal2 s 55272 0 55328 400 6 la_oenb[66]
port 462 nsew signal input
rlabel metal2 s 55776 0 55832 400 6 la_oenb[67]
port 463 nsew signal input
rlabel metal2 s 56280 0 56336 400 6 la_oenb[68]
port 464 nsew signal input
rlabel metal2 s 56784 0 56840 400 6 la_oenb[69]
port 465 nsew signal input
rlabel metal2 s 25032 0 25088 400 6 la_oenb[6]
port 466 nsew signal input
rlabel metal2 s 57288 0 57344 400 6 la_oenb[70]
port 467 nsew signal input
rlabel metal2 s 57792 0 57848 400 6 la_oenb[71]
port 468 nsew signal input
rlabel metal2 s 58296 0 58352 400 6 la_oenb[72]
port 469 nsew signal input
rlabel metal2 s 58800 0 58856 400 6 la_oenb[73]
port 470 nsew signal input
rlabel metal2 s 59304 0 59360 400 6 la_oenb[74]
port 471 nsew signal input
rlabel metal2 s 59808 0 59864 400 6 la_oenb[75]
port 472 nsew signal input
rlabel metal2 s 60312 0 60368 400 6 la_oenb[76]
port 473 nsew signal input
rlabel metal2 s 60816 0 60872 400 6 la_oenb[77]
port 474 nsew signal input
rlabel metal2 s 61320 0 61376 400 6 la_oenb[78]
port 475 nsew signal input
rlabel metal2 s 61824 0 61880 400 6 la_oenb[79]
port 476 nsew signal input
rlabel metal2 s 25536 0 25592 400 6 la_oenb[7]
port 477 nsew signal input
rlabel metal2 s 62328 0 62384 400 6 la_oenb[80]
port 478 nsew signal input
rlabel metal2 s 62832 0 62888 400 6 la_oenb[81]
port 479 nsew signal input
rlabel metal2 s 63336 0 63392 400 6 la_oenb[82]
port 480 nsew signal input
rlabel metal2 s 63840 0 63896 400 6 la_oenb[83]
port 481 nsew signal input
rlabel metal2 s 64344 0 64400 400 6 la_oenb[84]
port 482 nsew signal input
rlabel metal2 s 64848 0 64904 400 6 la_oenb[85]
port 483 nsew signal input
rlabel metal2 s 65352 0 65408 400 6 la_oenb[86]
port 484 nsew signal input
rlabel metal2 s 65856 0 65912 400 6 la_oenb[87]
port 485 nsew signal input
rlabel metal2 s 66360 0 66416 400 6 la_oenb[88]
port 486 nsew signal input
rlabel metal2 s 66864 0 66920 400 6 la_oenb[89]
port 487 nsew signal input
rlabel metal2 s 26040 0 26096 400 6 la_oenb[8]
port 488 nsew signal input
rlabel metal2 s 67368 0 67424 400 6 la_oenb[90]
port 489 nsew signal input
rlabel metal2 s 67872 0 67928 400 6 la_oenb[91]
port 490 nsew signal input
rlabel metal2 s 68376 0 68432 400 6 la_oenb[92]
port 491 nsew signal input
rlabel metal2 s 68880 0 68936 400 6 la_oenb[93]
port 492 nsew signal input
rlabel metal2 s 69384 0 69440 400 6 la_oenb[94]
port 493 nsew signal input
rlabel metal2 s 69888 0 69944 400 6 la_oenb[95]
port 494 nsew signal input
rlabel metal2 s 70392 0 70448 400 6 la_oenb[96]
port 495 nsew signal input
rlabel metal2 s 70896 0 70952 400 6 la_oenb[97]
port 496 nsew signal input
rlabel metal2 s 71400 0 71456 400 6 la_oenb[98]
port 497 nsew signal input
rlabel metal2 s 71904 0 71960 400 6 la_oenb[99]
port 498 nsew signal input
rlabel metal2 s 26544 0 26600 400 6 la_oenb[9]
port 499 nsew signal input
rlabel metal4 s 2224 1538 2384 58438 6 vdd
port 500 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 58438 6 vdd
port 500 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 58438 6 vdd
port 500 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 58438 6 vdd
port 500 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 58438 6 vdd
port 500 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 58438 6 vdd
port 500 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 58438 6 vss
port 501 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 58438 6 vss
port 501 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 58438 6 vss
port 501 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 58438 6 vss
port 501 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 58438 6 vss
port 501 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 58438 6 vss
port 501 nsew ground bidirectional
rlabel metal2 s 3864 0 3920 400 6 wb_clk_i
port 502 nsew signal input
rlabel metal2 s 4032 0 4088 400 6 wb_rst_i
port 503 nsew signal input
rlabel metal2 s 4200 0 4256 400 6 wbs_ack_o
port 504 nsew signal output
rlabel metal2 s 4872 0 4928 400 6 wbs_adr_i[0]
port 505 nsew signal input
rlabel metal2 s 10584 0 10640 400 6 wbs_adr_i[10]
port 506 nsew signal input
rlabel metal2 s 11088 0 11144 400 6 wbs_adr_i[11]
port 507 nsew signal input
rlabel metal2 s 11592 0 11648 400 6 wbs_adr_i[12]
port 508 nsew signal input
rlabel metal2 s 12096 0 12152 400 6 wbs_adr_i[13]
port 509 nsew signal input
rlabel metal2 s 12600 0 12656 400 6 wbs_adr_i[14]
port 510 nsew signal input
rlabel metal2 s 13104 0 13160 400 6 wbs_adr_i[15]
port 511 nsew signal input
rlabel metal2 s 13608 0 13664 400 6 wbs_adr_i[16]
port 512 nsew signal input
rlabel metal2 s 14112 0 14168 400 6 wbs_adr_i[17]
port 513 nsew signal input
rlabel metal2 s 14616 0 14672 400 6 wbs_adr_i[18]
port 514 nsew signal input
rlabel metal2 s 15120 0 15176 400 6 wbs_adr_i[19]
port 515 nsew signal input
rlabel metal2 s 5544 0 5600 400 6 wbs_adr_i[1]
port 516 nsew signal input
rlabel metal2 s 15624 0 15680 400 6 wbs_adr_i[20]
port 517 nsew signal input
rlabel metal2 s 16128 0 16184 400 6 wbs_adr_i[21]
port 518 nsew signal input
rlabel metal2 s 16632 0 16688 400 6 wbs_adr_i[22]
port 519 nsew signal input
rlabel metal2 s 17136 0 17192 400 6 wbs_adr_i[23]
port 520 nsew signal input
rlabel metal2 s 17640 0 17696 400 6 wbs_adr_i[24]
port 521 nsew signal input
rlabel metal2 s 18144 0 18200 400 6 wbs_adr_i[25]
port 522 nsew signal input
rlabel metal2 s 18648 0 18704 400 6 wbs_adr_i[26]
port 523 nsew signal input
rlabel metal2 s 19152 0 19208 400 6 wbs_adr_i[27]
port 524 nsew signal input
rlabel metal2 s 19656 0 19712 400 6 wbs_adr_i[28]
port 525 nsew signal input
rlabel metal2 s 20160 0 20216 400 6 wbs_adr_i[29]
port 526 nsew signal input
rlabel metal2 s 6216 0 6272 400 6 wbs_adr_i[2]
port 527 nsew signal input
rlabel metal2 s 20664 0 20720 400 6 wbs_adr_i[30]
port 528 nsew signal input
rlabel metal2 s 21168 0 21224 400 6 wbs_adr_i[31]
port 529 nsew signal input
rlabel metal2 s 6888 0 6944 400 6 wbs_adr_i[3]
port 530 nsew signal input
rlabel metal2 s 7560 0 7616 400 6 wbs_adr_i[4]
port 531 nsew signal input
rlabel metal2 s 8064 0 8120 400 6 wbs_adr_i[5]
port 532 nsew signal input
rlabel metal2 s 8568 0 8624 400 6 wbs_adr_i[6]
port 533 nsew signal input
rlabel metal2 s 9072 0 9128 400 6 wbs_adr_i[7]
port 534 nsew signal input
rlabel metal2 s 9576 0 9632 400 6 wbs_adr_i[8]
port 535 nsew signal input
rlabel metal2 s 10080 0 10136 400 6 wbs_adr_i[9]
port 536 nsew signal input
rlabel metal2 s 4368 0 4424 400 6 wbs_cyc_i
port 537 nsew signal input
rlabel metal2 s 5040 0 5096 400 6 wbs_dat_i[0]
port 538 nsew signal input
rlabel metal2 s 10752 0 10808 400 6 wbs_dat_i[10]
port 539 nsew signal input
rlabel metal2 s 11256 0 11312 400 6 wbs_dat_i[11]
port 540 nsew signal input
rlabel metal2 s 11760 0 11816 400 6 wbs_dat_i[12]
port 541 nsew signal input
rlabel metal2 s 12264 0 12320 400 6 wbs_dat_i[13]
port 542 nsew signal input
rlabel metal2 s 12768 0 12824 400 6 wbs_dat_i[14]
port 543 nsew signal input
rlabel metal2 s 13272 0 13328 400 6 wbs_dat_i[15]
port 544 nsew signal input
rlabel metal2 s 13776 0 13832 400 6 wbs_dat_i[16]
port 545 nsew signal input
rlabel metal2 s 14280 0 14336 400 6 wbs_dat_i[17]
port 546 nsew signal input
rlabel metal2 s 14784 0 14840 400 6 wbs_dat_i[18]
port 547 nsew signal input
rlabel metal2 s 15288 0 15344 400 6 wbs_dat_i[19]
port 548 nsew signal input
rlabel metal2 s 5712 0 5768 400 6 wbs_dat_i[1]
port 549 nsew signal input
rlabel metal2 s 15792 0 15848 400 6 wbs_dat_i[20]
port 550 nsew signal input
rlabel metal2 s 16296 0 16352 400 6 wbs_dat_i[21]
port 551 nsew signal input
rlabel metal2 s 16800 0 16856 400 6 wbs_dat_i[22]
port 552 nsew signal input
rlabel metal2 s 17304 0 17360 400 6 wbs_dat_i[23]
port 553 nsew signal input
rlabel metal2 s 17808 0 17864 400 6 wbs_dat_i[24]
port 554 nsew signal input
rlabel metal2 s 18312 0 18368 400 6 wbs_dat_i[25]
port 555 nsew signal input
rlabel metal2 s 18816 0 18872 400 6 wbs_dat_i[26]
port 556 nsew signal input
rlabel metal2 s 19320 0 19376 400 6 wbs_dat_i[27]
port 557 nsew signal input
rlabel metal2 s 19824 0 19880 400 6 wbs_dat_i[28]
port 558 nsew signal input
rlabel metal2 s 20328 0 20384 400 6 wbs_dat_i[29]
port 559 nsew signal input
rlabel metal2 s 6384 0 6440 400 6 wbs_dat_i[2]
port 560 nsew signal input
rlabel metal2 s 20832 0 20888 400 6 wbs_dat_i[30]
port 561 nsew signal input
rlabel metal2 s 21336 0 21392 400 6 wbs_dat_i[31]
port 562 nsew signal input
rlabel metal2 s 7056 0 7112 400 6 wbs_dat_i[3]
port 563 nsew signal input
rlabel metal2 s 7728 0 7784 400 6 wbs_dat_i[4]
port 564 nsew signal input
rlabel metal2 s 8232 0 8288 400 6 wbs_dat_i[5]
port 565 nsew signal input
rlabel metal2 s 8736 0 8792 400 6 wbs_dat_i[6]
port 566 nsew signal input
rlabel metal2 s 9240 0 9296 400 6 wbs_dat_i[7]
port 567 nsew signal input
rlabel metal2 s 9744 0 9800 400 6 wbs_dat_i[8]
port 568 nsew signal input
rlabel metal2 s 10248 0 10304 400 6 wbs_dat_i[9]
port 569 nsew signal input
rlabel metal2 s 5208 0 5264 400 6 wbs_dat_o[0]
port 570 nsew signal output
rlabel metal2 s 10920 0 10976 400 6 wbs_dat_o[10]
port 571 nsew signal output
rlabel metal2 s 11424 0 11480 400 6 wbs_dat_o[11]
port 572 nsew signal output
rlabel metal2 s 11928 0 11984 400 6 wbs_dat_o[12]
port 573 nsew signal output
rlabel metal2 s 12432 0 12488 400 6 wbs_dat_o[13]
port 574 nsew signal output
rlabel metal2 s 12936 0 12992 400 6 wbs_dat_o[14]
port 575 nsew signal output
rlabel metal2 s 13440 0 13496 400 6 wbs_dat_o[15]
port 576 nsew signal output
rlabel metal2 s 13944 0 14000 400 6 wbs_dat_o[16]
port 577 nsew signal output
rlabel metal2 s 14448 0 14504 400 6 wbs_dat_o[17]
port 578 nsew signal output
rlabel metal2 s 14952 0 15008 400 6 wbs_dat_o[18]
port 579 nsew signal output
rlabel metal2 s 15456 0 15512 400 6 wbs_dat_o[19]
port 580 nsew signal output
rlabel metal2 s 5880 0 5936 400 6 wbs_dat_o[1]
port 581 nsew signal output
rlabel metal2 s 15960 0 16016 400 6 wbs_dat_o[20]
port 582 nsew signal output
rlabel metal2 s 16464 0 16520 400 6 wbs_dat_o[21]
port 583 nsew signal output
rlabel metal2 s 16968 0 17024 400 6 wbs_dat_o[22]
port 584 nsew signal output
rlabel metal2 s 17472 0 17528 400 6 wbs_dat_o[23]
port 585 nsew signal output
rlabel metal2 s 17976 0 18032 400 6 wbs_dat_o[24]
port 586 nsew signal output
rlabel metal2 s 18480 0 18536 400 6 wbs_dat_o[25]
port 587 nsew signal output
rlabel metal2 s 18984 0 19040 400 6 wbs_dat_o[26]
port 588 nsew signal output
rlabel metal2 s 19488 0 19544 400 6 wbs_dat_o[27]
port 589 nsew signal output
rlabel metal2 s 19992 0 20048 400 6 wbs_dat_o[28]
port 590 nsew signal output
rlabel metal2 s 20496 0 20552 400 6 wbs_dat_o[29]
port 591 nsew signal output
rlabel metal2 s 6552 0 6608 400 6 wbs_dat_o[2]
port 592 nsew signal output
rlabel metal2 s 21000 0 21056 400 6 wbs_dat_o[30]
port 593 nsew signal output
rlabel metal2 s 21504 0 21560 400 6 wbs_dat_o[31]
port 594 nsew signal output
rlabel metal2 s 7224 0 7280 400 6 wbs_dat_o[3]
port 595 nsew signal output
rlabel metal2 s 7896 0 7952 400 6 wbs_dat_o[4]
port 596 nsew signal output
rlabel metal2 s 8400 0 8456 400 6 wbs_dat_o[5]
port 597 nsew signal output
rlabel metal2 s 8904 0 8960 400 6 wbs_dat_o[6]
port 598 nsew signal output
rlabel metal2 s 9408 0 9464 400 6 wbs_dat_o[7]
port 599 nsew signal output
rlabel metal2 s 9912 0 9968 400 6 wbs_dat_o[8]
port 600 nsew signal output
rlabel metal2 s 10416 0 10472 400 6 wbs_dat_o[9]
port 601 nsew signal output
rlabel metal2 s 5376 0 5432 400 6 wbs_sel_i[0]
port 602 nsew signal input
rlabel metal2 s 6048 0 6104 400 6 wbs_sel_i[1]
port 603 nsew signal input
rlabel metal2 s 6720 0 6776 400 6 wbs_sel_i[2]
port 604 nsew signal input
rlabel metal2 s 7392 0 7448 400 6 wbs_sel_i[3]
port 605 nsew signal input
rlabel metal2 s 4536 0 4592 400 6 wbs_stb_i
port 606 nsew signal input
rlabel metal2 s 4704 0 4760 400 6 wbs_we_i
port 607 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 90000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2526888
string GDS_FILE /opt/caravel_180/openlane/user_proj_example/runs/22_12_03_04_01/results/signoff/macro_golden.magic.gds
string GDS_START 169586
<< end >>

