magic
tech gf180mcuC
magscale 1 5
timestamp 1670243369
<< obsm1 >>
rect 118172 169855 176804 231153
<< metal2 >>
rect 4900 297780 5012 298500
rect 13132 297780 13244 298500
rect 21364 297780 21476 298500
rect 29596 297780 29708 298500
rect 37828 297780 37940 298500
rect 46060 297780 46172 298500
rect 54292 297780 54404 298500
rect 62524 297780 62636 298500
rect 70756 297780 70868 298500
rect 78988 297780 79100 298500
rect 87220 297780 87332 298500
rect 95452 297780 95564 298500
rect 103684 297780 103796 298500
rect 111916 297780 112028 298500
rect 120148 297780 120260 298500
rect 128380 297780 128492 298500
rect 136612 297780 136724 298500
rect 144844 297780 144956 298500
rect 153076 297780 153188 298500
rect 161308 297780 161420 298500
rect 169540 297780 169652 298500
rect 177772 297780 177884 298500
rect 186004 297780 186116 298500
rect 194236 297780 194348 298500
rect 202468 297780 202580 298500
rect 210700 297780 210812 298500
rect 218932 297780 219044 298500
rect 227164 297780 227276 298500
rect 235396 297780 235508 298500
rect 243628 297780 243740 298500
rect 251860 297780 251972 298500
rect 260092 297780 260204 298500
rect 268324 297780 268436 298500
rect 276556 297780 276668 298500
rect 284788 297780 284900 298500
rect 293020 297780 293132 298500
rect 5684 -480 5796 240
rect 6636 -480 6748 240
rect 7588 -480 7700 240
rect 8540 -480 8652 240
rect 9492 -480 9604 240
rect 10444 -480 10556 240
rect 11396 -480 11508 240
rect 12348 -480 12460 240
rect 13300 -480 13412 240
rect 14252 -480 14364 240
rect 15204 -480 15316 240
rect 16156 -480 16268 240
rect 17108 -480 17220 240
rect 18060 -480 18172 240
rect 19012 -480 19124 240
rect 19964 -480 20076 240
rect 20916 -480 21028 240
rect 21868 -480 21980 240
rect 22820 -480 22932 240
rect 23772 -480 23884 240
rect 24724 -480 24836 240
rect 25676 -480 25788 240
rect 26628 -480 26740 240
rect 27580 -480 27692 240
rect 28532 -480 28644 240
rect 29484 -480 29596 240
rect 30436 -480 30548 240
rect 31388 -480 31500 240
rect 32340 -480 32452 240
rect 33292 -480 33404 240
rect 34244 -480 34356 240
rect 35196 -480 35308 240
rect 36148 -480 36260 240
rect 37100 -480 37212 240
rect 38052 -480 38164 240
rect 39004 -480 39116 240
rect 39956 -480 40068 240
rect 40908 -480 41020 240
rect 41860 -480 41972 240
rect 42812 -480 42924 240
rect 43764 -480 43876 240
rect 44716 -480 44828 240
rect 45668 -480 45780 240
rect 46620 -480 46732 240
rect 47572 -480 47684 240
rect 48524 -480 48636 240
rect 49476 -480 49588 240
rect 50428 -480 50540 240
rect 51380 -480 51492 240
rect 52332 -480 52444 240
rect 53284 -480 53396 240
rect 54236 -480 54348 240
rect 55188 -480 55300 240
rect 56140 -480 56252 240
rect 57092 -480 57204 240
rect 58044 -480 58156 240
rect 58996 -480 59108 240
rect 59948 -480 60060 240
rect 60900 -480 61012 240
rect 61852 -480 61964 240
rect 62804 -480 62916 240
rect 63756 -480 63868 240
rect 64708 -480 64820 240
rect 65660 -480 65772 240
rect 66612 -480 66724 240
rect 67564 -480 67676 240
rect 68516 -480 68628 240
rect 69468 -480 69580 240
rect 70420 -480 70532 240
rect 71372 -480 71484 240
rect 72324 -480 72436 240
rect 73276 -480 73388 240
rect 74228 -480 74340 240
rect 75180 -480 75292 240
rect 76132 -480 76244 240
rect 77084 -480 77196 240
rect 78036 -480 78148 240
rect 78988 -480 79100 240
rect 79940 -480 80052 240
rect 80892 -480 81004 240
rect 81844 -480 81956 240
rect 82796 -480 82908 240
rect 83748 -480 83860 240
rect 84700 -480 84812 240
rect 85652 -480 85764 240
rect 86604 -480 86716 240
rect 87556 -480 87668 240
rect 88508 -480 88620 240
rect 89460 -480 89572 240
rect 90412 -480 90524 240
rect 91364 -480 91476 240
rect 92316 -480 92428 240
rect 93268 -480 93380 240
rect 94220 -480 94332 240
rect 95172 -480 95284 240
rect 96124 -480 96236 240
rect 97076 -480 97188 240
rect 98028 -480 98140 240
rect 98980 -480 99092 240
rect 99932 -480 100044 240
rect 100884 -480 100996 240
rect 101836 -480 101948 240
rect 102788 -480 102900 240
rect 103740 -480 103852 240
rect 104692 -480 104804 240
rect 105644 -480 105756 240
rect 106596 -480 106708 240
rect 107548 -480 107660 240
rect 108500 -480 108612 240
rect 109452 -480 109564 240
rect 110404 -480 110516 240
rect 111356 -480 111468 240
rect 112308 -480 112420 240
rect 113260 -480 113372 240
rect 114212 -480 114324 240
rect 115164 -480 115276 240
rect 116116 -480 116228 240
rect 117068 -480 117180 240
rect 118020 -480 118132 240
rect 118972 -480 119084 240
rect 119924 -480 120036 240
rect 120876 -480 120988 240
rect 121828 -480 121940 240
rect 122780 -480 122892 240
rect 123732 -480 123844 240
rect 124684 -480 124796 240
rect 125636 -480 125748 240
rect 126588 -480 126700 240
rect 127540 -480 127652 240
rect 128492 -480 128604 240
rect 129444 -480 129556 240
rect 130396 -480 130508 240
rect 131348 -480 131460 240
rect 132300 -480 132412 240
rect 133252 -480 133364 240
rect 134204 -480 134316 240
rect 135156 -480 135268 240
rect 136108 -480 136220 240
rect 137060 -480 137172 240
rect 138012 -480 138124 240
rect 138964 -480 139076 240
rect 139916 -480 140028 240
rect 140868 -480 140980 240
rect 141820 -480 141932 240
rect 142772 -480 142884 240
rect 143724 -480 143836 240
rect 144676 -480 144788 240
rect 145628 -480 145740 240
rect 146580 -480 146692 240
rect 147532 -480 147644 240
rect 148484 -480 148596 240
rect 149436 -480 149548 240
rect 150388 -480 150500 240
rect 151340 -480 151452 240
rect 152292 -480 152404 240
rect 153244 -480 153356 240
rect 154196 -480 154308 240
rect 155148 -480 155260 240
rect 156100 -480 156212 240
rect 157052 -480 157164 240
rect 158004 -480 158116 240
rect 158956 -480 159068 240
rect 159908 -480 160020 240
rect 160860 -480 160972 240
rect 161812 -480 161924 240
rect 162764 -480 162876 240
rect 163716 -480 163828 240
rect 164668 -480 164780 240
rect 165620 -480 165732 240
rect 166572 -480 166684 240
rect 167524 -480 167636 240
rect 168476 -480 168588 240
rect 169428 -480 169540 240
rect 170380 -480 170492 240
rect 171332 -480 171444 240
rect 172284 -480 172396 240
rect 173236 -480 173348 240
rect 174188 -480 174300 240
rect 175140 -480 175252 240
rect 176092 -480 176204 240
rect 177044 -480 177156 240
rect 177996 -480 178108 240
rect 178948 -480 179060 240
rect 179900 -480 180012 240
rect 180852 -480 180964 240
rect 181804 -480 181916 240
rect 182756 -480 182868 240
rect 183708 -480 183820 240
rect 184660 -480 184772 240
rect 185612 -480 185724 240
rect 186564 -480 186676 240
rect 187516 -480 187628 240
rect 188468 -480 188580 240
rect 189420 -480 189532 240
rect 190372 -480 190484 240
rect 191324 -480 191436 240
rect 192276 -480 192388 240
rect 193228 -480 193340 240
rect 194180 -480 194292 240
rect 195132 -480 195244 240
rect 196084 -480 196196 240
rect 197036 -480 197148 240
rect 197988 -480 198100 240
rect 198940 -480 199052 240
rect 199892 -480 200004 240
rect 200844 -480 200956 240
rect 201796 -480 201908 240
rect 202748 -480 202860 240
rect 203700 -480 203812 240
rect 204652 -480 204764 240
rect 205604 -480 205716 240
rect 206556 -480 206668 240
rect 207508 -480 207620 240
rect 208460 -480 208572 240
rect 209412 -480 209524 240
rect 210364 -480 210476 240
rect 211316 -480 211428 240
rect 212268 -480 212380 240
rect 213220 -480 213332 240
rect 214172 -480 214284 240
rect 215124 -480 215236 240
rect 216076 -480 216188 240
rect 217028 -480 217140 240
rect 217980 -480 218092 240
rect 218932 -480 219044 240
rect 219884 -480 219996 240
rect 220836 -480 220948 240
rect 221788 -480 221900 240
rect 222740 -480 222852 240
rect 223692 -480 223804 240
rect 224644 -480 224756 240
rect 225596 -480 225708 240
rect 226548 -480 226660 240
rect 227500 -480 227612 240
rect 228452 -480 228564 240
rect 229404 -480 229516 240
rect 230356 -480 230468 240
rect 231308 -480 231420 240
rect 232260 -480 232372 240
rect 233212 -480 233324 240
rect 234164 -480 234276 240
rect 235116 -480 235228 240
rect 236068 -480 236180 240
rect 237020 -480 237132 240
rect 237972 -480 238084 240
rect 238924 -480 239036 240
rect 239876 -480 239988 240
rect 240828 -480 240940 240
rect 241780 -480 241892 240
rect 242732 -480 242844 240
rect 243684 -480 243796 240
rect 244636 -480 244748 240
rect 245588 -480 245700 240
rect 246540 -480 246652 240
rect 247492 -480 247604 240
rect 248444 -480 248556 240
rect 249396 -480 249508 240
rect 250348 -480 250460 240
rect 251300 -480 251412 240
rect 252252 -480 252364 240
rect 253204 -480 253316 240
rect 254156 -480 254268 240
rect 255108 -480 255220 240
rect 256060 -480 256172 240
rect 257012 -480 257124 240
rect 257964 -480 258076 240
rect 258916 -480 259028 240
rect 259868 -480 259980 240
rect 260820 -480 260932 240
rect 261772 -480 261884 240
rect 262724 -480 262836 240
rect 263676 -480 263788 240
rect 264628 -480 264740 240
rect 265580 -480 265692 240
rect 266532 -480 266644 240
rect 267484 -480 267596 240
rect 268436 -480 268548 240
rect 269388 -480 269500 240
rect 270340 -480 270452 240
rect 271292 -480 271404 240
rect 272244 -480 272356 240
rect 273196 -480 273308 240
rect 274148 -480 274260 240
rect 275100 -480 275212 240
rect 276052 -480 276164 240
rect 277004 -480 277116 240
rect 277956 -480 278068 240
rect 278908 -480 279020 240
rect 279860 -480 279972 240
rect 280812 -480 280924 240
rect 281764 -480 281876 240
rect 282716 -480 282828 240
rect 283668 -480 283780 240
rect 284620 -480 284732 240
rect 285572 -480 285684 240
rect 286524 -480 286636 240
rect 287476 -480 287588 240
rect 288428 -480 288540 240
rect 289380 -480 289492 240
rect 290332 -480 290444 240
rect 291284 -480 291396 240
rect 292236 -480 292348 240
<< obsm2 >>
rect 2926 297750 4870 297850
rect 5042 297750 13102 297850
rect 13274 297750 21334 297850
rect 21506 297750 29566 297850
rect 29738 297750 37798 297850
rect 37970 297750 46030 297850
rect 46202 297750 54262 297850
rect 54434 297750 62494 297850
rect 62666 297750 70726 297850
rect 70898 297750 78958 297850
rect 79130 297750 87190 297850
rect 87362 297750 95422 297850
rect 95594 297750 103654 297850
rect 103826 297750 111886 297850
rect 112058 297750 120118 297850
rect 120290 297750 128350 297850
rect 128522 297750 136582 297850
rect 136754 297750 144814 297850
rect 144986 297750 153046 297850
rect 153218 297750 161278 297850
rect 161450 297750 169510 297850
rect 169682 297750 177742 297850
rect 177914 297750 185974 297850
rect 186146 297750 194206 297850
rect 194378 297750 202438 297850
rect 202610 297750 210670 297850
rect 210842 297750 218902 297850
rect 219074 297750 227134 297850
rect 227306 297750 235366 297850
rect 235538 297750 243598 297850
rect 243770 297750 251830 297850
rect 252002 297750 260062 297850
rect 260234 297750 268294 297850
rect 268466 297750 276526 297850
rect 276698 297750 284758 297850
rect 284930 297750 292990 297850
rect 293162 297750 297010 297850
rect 2926 270 297010 297750
rect 2926 182 5654 270
rect 5826 182 6606 270
rect 6778 182 7558 270
rect 7730 182 8510 270
rect 8682 182 9462 270
rect 9634 182 10414 270
rect 10586 182 11366 270
rect 11538 182 12318 270
rect 12490 182 13270 270
rect 13442 182 14222 270
rect 14394 182 15174 270
rect 15346 182 16126 270
rect 16298 182 17078 270
rect 17250 182 18030 270
rect 18202 182 18982 270
rect 19154 182 19934 270
rect 20106 182 20886 270
rect 21058 182 21838 270
rect 22010 182 22790 270
rect 22962 182 23742 270
rect 23914 182 24694 270
rect 24866 182 25646 270
rect 25818 182 26598 270
rect 26770 182 27550 270
rect 27722 182 28502 270
rect 28674 182 29454 270
rect 29626 182 30406 270
rect 30578 182 31358 270
rect 31530 182 32310 270
rect 32482 182 33262 270
rect 33434 182 34214 270
rect 34386 182 35166 270
rect 35338 182 36118 270
rect 36290 182 37070 270
rect 37242 182 38022 270
rect 38194 182 38974 270
rect 39146 182 39926 270
rect 40098 182 40878 270
rect 41050 182 41830 270
rect 42002 182 42782 270
rect 42954 182 43734 270
rect 43906 182 44686 270
rect 44858 182 45638 270
rect 45810 182 46590 270
rect 46762 182 47542 270
rect 47714 182 48494 270
rect 48666 182 49446 270
rect 49618 182 50398 270
rect 50570 182 51350 270
rect 51522 182 52302 270
rect 52474 182 53254 270
rect 53426 182 54206 270
rect 54378 182 55158 270
rect 55330 182 56110 270
rect 56282 182 57062 270
rect 57234 182 58014 270
rect 58186 182 58966 270
rect 59138 182 59918 270
rect 60090 182 60870 270
rect 61042 182 61822 270
rect 61994 182 62774 270
rect 62946 182 63726 270
rect 63898 182 64678 270
rect 64850 182 65630 270
rect 65802 182 66582 270
rect 66754 182 67534 270
rect 67706 182 68486 270
rect 68658 182 69438 270
rect 69610 182 70390 270
rect 70562 182 71342 270
rect 71514 182 72294 270
rect 72466 182 73246 270
rect 73418 182 74198 270
rect 74370 182 75150 270
rect 75322 182 76102 270
rect 76274 182 77054 270
rect 77226 182 78006 270
rect 78178 182 78958 270
rect 79130 182 79910 270
rect 80082 182 80862 270
rect 81034 182 81814 270
rect 81986 182 82766 270
rect 82938 182 83718 270
rect 83890 182 84670 270
rect 84842 182 85622 270
rect 85794 182 86574 270
rect 86746 182 87526 270
rect 87698 182 88478 270
rect 88650 182 89430 270
rect 89602 182 90382 270
rect 90554 182 91334 270
rect 91506 182 92286 270
rect 92458 182 93238 270
rect 93410 182 94190 270
rect 94362 182 95142 270
rect 95314 182 96094 270
rect 96266 182 97046 270
rect 97218 182 97998 270
rect 98170 182 98950 270
rect 99122 182 99902 270
rect 100074 182 100854 270
rect 101026 182 101806 270
rect 101978 182 102758 270
rect 102930 182 103710 270
rect 103882 182 104662 270
rect 104834 182 105614 270
rect 105786 182 106566 270
rect 106738 182 107518 270
rect 107690 182 108470 270
rect 108642 182 109422 270
rect 109594 182 110374 270
rect 110546 182 111326 270
rect 111498 182 112278 270
rect 112450 182 113230 270
rect 113402 182 114182 270
rect 114354 182 115134 270
rect 115306 182 116086 270
rect 116258 182 117038 270
rect 117210 182 117990 270
rect 118162 182 118942 270
rect 119114 182 119894 270
rect 120066 182 120846 270
rect 121018 182 121798 270
rect 121970 182 122750 270
rect 122922 182 123702 270
rect 123874 182 124654 270
rect 124826 182 125606 270
rect 125778 182 126558 270
rect 126730 182 127510 270
rect 127682 182 128462 270
rect 128634 182 129414 270
rect 129586 182 130366 270
rect 130538 182 131318 270
rect 131490 182 132270 270
rect 132442 182 133222 270
rect 133394 182 134174 270
rect 134346 182 135126 270
rect 135298 182 136078 270
rect 136250 182 137030 270
rect 137202 182 137982 270
rect 138154 182 138934 270
rect 139106 182 139886 270
rect 140058 182 140838 270
rect 141010 182 141790 270
rect 141962 182 142742 270
rect 142914 182 143694 270
rect 143866 182 144646 270
rect 144818 182 145598 270
rect 145770 182 146550 270
rect 146722 182 147502 270
rect 147674 182 148454 270
rect 148626 182 149406 270
rect 149578 182 150358 270
rect 150530 182 151310 270
rect 151482 182 152262 270
rect 152434 182 153214 270
rect 153386 182 154166 270
rect 154338 182 155118 270
rect 155290 182 156070 270
rect 156242 182 157022 270
rect 157194 182 157974 270
rect 158146 182 158926 270
rect 159098 182 159878 270
rect 160050 182 160830 270
rect 161002 182 161782 270
rect 161954 182 162734 270
rect 162906 182 163686 270
rect 163858 182 164638 270
rect 164810 182 165590 270
rect 165762 182 166542 270
rect 166714 182 167494 270
rect 167666 182 168446 270
rect 168618 182 169398 270
rect 169570 182 170350 270
rect 170522 182 171302 270
rect 171474 182 172254 270
rect 172426 182 173206 270
rect 173378 182 174158 270
rect 174330 182 175110 270
rect 175282 182 176062 270
rect 176234 182 177014 270
rect 177186 182 177966 270
rect 178138 182 178918 270
rect 179090 182 179870 270
rect 180042 182 180822 270
rect 180994 182 181774 270
rect 181946 182 182726 270
rect 182898 182 183678 270
rect 183850 182 184630 270
rect 184802 182 185582 270
rect 185754 182 186534 270
rect 186706 182 187486 270
rect 187658 182 188438 270
rect 188610 182 189390 270
rect 189562 182 190342 270
rect 190514 182 191294 270
rect 191466 182 192246 270
rect 192418 182 193198 270
rect 193370 182 194150 270
rect 194322 182 195102 270
rect 195274 182 196054 270
rect 196226 182 197006 270
rect 197178 182 197958 270
rect 198130 182 198910 270
rect 199082 182 199862 270
rect 200034 182 200814 270
rect 200986 182 201766 270
rect 201938 182 202718 270
rect 202890 182 203670 270
rect 203842 182 204622 270
rect 204794 182 205574 270
rect 205746 182 206526 270
rect 206698 182 207478 270
rect 207650 182 208430 270
rect 208602 182 209382 270
rect 209554 182 210334 270
rect 210506 182 211286 270
rect 211458 182 212238 270
rect 212410 182 213190 270
rect 213362 182 214142 270
rect 214314 182 215094 270
rect 215266 182 216046 270
rect 216218 182 216998 270
rect 217170 182 217950 270
rect 218122 182 218902 270
rect 219074 182 219854 270
rect 220026 182 220806 270
rect 220978 182 221758 270
rect 221930 182 222710 270
rect 222882 182 223662 270
rect 223834 182 224614 270
rect 224786 182 225566 270
rect 225738 182 226518 270
rect 226690 182 227470 270
rect 227642 182 228422 270
rect 228594 182 229374 270
rect 229546 182 230326 270
rect 230498 182 231278 270
rect 231450 182 232230 270
rect 232402 182 233182 270
rect 233354 182 234134 270
rect 234306 182 235086 270
rect 235258 182 236038 270
rect 236210 182 236990 270
rect 237162 182 237942 270
rect 238114 182 238894 270
rect 239066 182 239846 270
rect 240018 182 240798 270
rect 240970 182 241750 270
rect 241922 182 242702 270
rect 242874 182 243654 270
rect 243826 182 244606 270
rect 244778 182 245558 270
rect 245730 182 246510 270
rect 246682 182 247462 270
rect 247634 182 248414 270
rect 248586 182 249366 270
rect 249538 182 250318 270
rect 250490 182 251270 270
rect 251442 182 252222 270
rect 252394 182 253174 270
rect 253346 182 254126 270
rect 254298 182 255078 270
rect 255250 182 256030 270
rect 256202 182 256982 270
rect 257154 182 257934 270
rect 258106 182 258886 270
rect 259058 182 259838 270
rect 260010 182 260790 270
rect 260962 182 261742 270
rect 261914 182 262694 270
rect 262866 182 263646 270
rect 263818 182 264598 270
rect 264770 182 265550 270
rect 265722 182 266502 270
rect 266674 182 267454 270
rect 267626 182 268406 270
rect 268578 182 269358 270
rect 269530 182 270310 270
rect 270482 182 271262 270
rect 271434 182 272214 270
rect 272386 182 273166 270
rect 273338 182 274118 270
rect 274290 182 275070 270
rect 275242 182 276022 270
rect 276194 182 276974 270
rect 277146 182 277926 270
rect 278098 182 278878 270
rect 279050 182 279830 270
rect 280002 182 280782 270
rect 280954 182 281734 270
rect 281906 182 282686 270
rect 282858 182 283638 270
rect 283810 182 284590 270
rect 284762 182 285542 270
rect 285714 182 286494 270
rect 286666 182 287446 270
rect 287618 182 288398 270
rect 288570 182 289350 270
rect 289522 182 290302 270
rect 290474 182 291254 270
rect 291426 182 292206 270
rect 292378 182 297010 270
<< metal3 >>
rect 297780 294532 298500 294644
rect -480 294364 240 294476
rect -480 288876 240 288988
rect 297780 288932 298500 289044
rect -480 283388 240 283500
rect 297780 283332 298500 283444
rect -480 277900 240 278012
rect 297780 277732 298500 277844
rect -480 272412 240 272524
rect 297780 272132 298500 272244
rect -480 266924 240 267036
rect 297780 266532 298500 266644
rect -480 261436 240 261548
rect 297780 260932 298500 261044
rect -480 255948 240 256060
rect 297780 255332 298500 255444
rect -480 250460 240 250572
rect 297780 249732 298500 249844
rect -480 244972 240 245084
rect 297780 244132 298500 244244
rect -480 239484 240 239596
rect 297780 238532 298500 238644
rect -480 233996 240 234108
rect 297780 232932 298500 233044
rect -480 228508 240 228620
rect 297780 227332 298500 227444
rect -480 223020 240 223132
rect 297780 221732 298500 221844
rect -480 217532 240 217644
rect 297780 216132 298500 216244
rect -480 212044 240 212156
rect 297780 210532 298500 210644
rect -480 206556 240 206668
rect 297780 204932 298500 205044
rect -480 201068 240 201180
rect 297780 199332 298500 199444
rect -480 195580 240 195692
rect 297780 193732 298500 193844
rect -480 190092 240 190204
rect 297780 188132 298500 188244
rect -480 184604 240 184716
rect 297780 182532 298500 182644
rect -480 179116 240 179228
rect 297780 176932 298500 177044
rect -480 173628 240 173740
rect 297780 171332 298500 171444
rect -480 168140 240 168252
rect 297780 165732 298500 165844
rect -480 162652 240 162764
rect 297780 160132 298500 160244
rect -480 157164 240 157276
rect 297780 154532 298500 154644
rect -480 151676 240 151788
rect 297780 148932 298500 149044
rect -480 146188 240 146300
rect 297780 143332 298500 143444
rect -480 140700 240 140812
rect 297780 137732 298500 137844
rect -480 135212 240 135324
rect 297780 132132 298500 132244
rect -480 129724 240 129836
rect 297780 126532 298500 126644
rect -480 124236 240 124348
rect 297780 120932 298500 121044
rect -480 118748 240 118860
rect 297780 115332 298500 115444
rect -480 113260 240 113372
rect 297780 109732 298500 109844
rect -480 107772 240 107884
rect 297780 104132 298500 104244
rect -480 102284 240 102396
rect 297780 98532 298500 98644
rect -480 96796 240 96908
rect 297780 92932 298500 93044
rect -480 91308 240 91420
rect 297780 87332 298500 87444
rect -480 85820 240 85932
rect 297780 81732 298500 81844
rect -480 80332 240 80444
rect 297780 76132 298500 76244
rect -480 74844 240 74956
rect 297780 70532 298500 70644
rect -480 69356 240 69468
rect 297780 64932 298500 65044
rect -480 63868 240 63980
rect 297780 59332 298500 59444
rect -480 58380 240 58492
rect 297780 53732 298500 53844
rect -480 52892 240 53004
rect 297780 48132 298500 48244
rect -480 47404 240 47516
rect 297780 42532 298500 42644
rect -480 41916 240 42028
rect 297780 36932 298500 37044
rect -480 36428 240 36540
rect 297780 31332 298500 31444
rect -480 30940 240 31052
rect 297780 25732 298500 25844
rect -480 25452 240 25564
rect 297780 20132 298500 20244
rect -480 19964 240 20076
rect -480 14476 240 14588
rect 297780 14532 298500 14644
rect -480 8988 240 9100
rect 297780 8932 298500 9044
rect -480 3500 240 3612
rect 297780 3332 298500 3444
<< obsm3 >>
rect 182 294674 297850 295666
rect 182 294506 297750 294674
rect 270 294502 297750 294506
rect 270 294334 297850 294502
rect 182 289074 297850 294334
rect 182 289018 297750 289074
rect 270 288902 297750 289018
rect 270 288846 297850 288902
rect 182 283530 297850 288846
rect 270 283474 297850 283530
rect 270 283358 297750 283474
rect 182 283302 297750 283358
rect 182 278042 297850 283302
rect 270 277874 297850 278042
rect 270 277870 297750 277874
rect 182 277702 297750 277870
rect 182 272554 297850 277702
rect 270 272382 297850 272554
rect 182 272274 297850 272382
rect 182 272102 297750 272274
rect 182 267066 297850 272102
rect 270 266894 297850 267066
rect 182 266674 297850 266894
rect 182 266502 297750 266674
rect 182 261578 297850 266502
rect 270 261406 297850 261578
rect 182 261074 297850 261406
rect 182 260902 297750 261074
rect 182 256090 297850 260902
rect 270 255918 297850 256090
rect 182 255474 297850 255918
rect 182 255302 297750 255474
rect 182 250602 297850 255302
rect 270 250430 297850 250602
rect 182 249874 297850 250430
rect 182 249702 297750 249874
rect 182 245114 297850 249702
rect 270 244942 297850 245114
rect 182 244274 297850 244942
rect 182 244102 297750 244274
rect 182 239626 297850 244102
rect 270 239454 297850 239626
rect 182 238674 297850 239454
rect 182 238502 297750 238674
rect 182 234138 297850 238502
rect 270 233966 297850 234138
rect 182 233074 297850 233966
rect 182 232902 297750 233074
rect 182 228650 297850 232902
rect 270 228478 297850 228650
rect 182 227474 297850 228478
rect 182 227302 297750 227474
rect 182 223162 297850 227302
rect 270 222990 297850 223162
rect 182 221874 297850 222990
rect 182 221702 297750 221874
rect 182 217674 297850 221702
rect 270 217502 297850 217674
rect 182 216274 297850 217502
rect 182 216102 297750 216274
rect 182 212186 297850 216102
rect 270 212014 297850 212186
rect 182 210674 297850 212014
rect 182 210502 297750 210674
rect 182 206698 297850 210502
rect 270 206526 297850 206698
rect 182 205074 297850 206526
rect 182 204902 297750 205074
rect 182 201210 297850 204902
rect 270 201038 297850 201210
rect 182 199474 297850 201038
rect 182 199302 297750 199474
rect 182 195722 297850 199302
rect 270 195550 297850 195722
rect 182 193874 297850 195550
rect 182 193702 297750 193874
rect 182 190234 297850 193702
rect 270 190062 297850 190234
rect 182 188274 297850 190062
rect 182 188102 297750 188274
rect 182 184746 297850 188102
rect 270 184574 297850 184746
rect 182 182674 297850 184574
rect 182 182502 297750 182674
rect 182 179258 297850 182502
rect 270 179086 297850 179258
rect 182 177074 297850 179086
rect 182 176902 297750 177074
rect 182 173770 297850 176902
rect 270 173598 297850 173770
rect 182 171474 297850 173598
rect 182 171302 297750 171474
rect 182 168282 297850 171302
rect 270 168110 297850 168282
rect 182 165874 297850 168110
rect 182 165702 297750 165874
rect 182 162794 297850 165702
rect 270 162622 297850 162794
rect 182 160274 297850 162622
rect 182 160102 297750 160274
rect 182 157306 297850 160102
rect 270 157134 297850 157306
rect 182 154674 297850 157134
rect 182 154502 297750 154674
rect 182 151818 297850 154502
rect 270 151646 297850 151818
rect 182 149074 297850 151646
rect 182 148902 297750 149074
rect 182 146330 297850 148902
rect 270 146158 297850 146330
rect 182 143474 297850 146158
rect 182 143302 297750 143474
rect 182 140842 297850 143302
rect 270 140670 297850 140842
rect 182 137874 297850 140670
rect 182 137702 297750 137874
rect 182 135354 297850 137702
rect 270 135182 297850 135354
rect 182 132274 297850 135182
rect 182 132102 297750 132274
rect 182 129866 297850 132102
rect 270 129694 297850 129866
rect 182 126674 297850 129694
rect 182 126502 297750 126674
rect 182 124378 297850 126502
rect 270 124206 297850 124378
rect 182 121074 297850 124206
rect 182 120902 297750 121074
rect 182 118890 297850 120902
rect 270 118718 297850 118890
rect 182 115474 297850 118718
rect 182 115302 297750 115474
rect 182 113402 297850 115302
rect 270 113230 297850 113402
rect 182 109874 297850 113230
rect 182 109702 297750 109874
rect 182 107914 297850 109702
rect 270 107742 297850 107914
rect 182 104274 297850 107742
rect 182 104102 297750 104274
rect 182 102426 297850 104102
rect 270 102254 297850 102426
rect 182 98674 297850 102254
rect 182 98502 297750 98674
rect 182 96938 297850 98502
rect 270 96766 297850 96938
rect 182 93074 297850 96766
rect 182 92902 297750 93074
rect 182 91450 297850 92902
rect 270 91278 297850 91450
rect 182 87474 297850 91278
rect 182 87302 297750 87474
rect 182 85962 297850 87302
rect 270 85790 297850 85962
rect 182 81874 297850 85790
rect 182 81702 297750 81874
rect 182 80474 297850 81702
rect 270 80302 297850 80474
rect 182 76274 297850 80302
rect 182 76102 297750 76274
rect 182 74986 297850 76102
rect 270 74814 297850 74986
rect 182 70674 297850 74814
rect 182 70502 297750 70674
rect 182 69498 297850 70502
rect 270 69326 297850 69498
rect 182 65074 297850 69326
rect 182 64902 297750 65074
rect 182 64010 297850 64902
rect 270 63838 297850 64010
rect 182 59474 297850 63838
rect 182 59302 297750 59474
rect 182 58522 297850 59302
rect 270 58350 297850 58522
rect 182 53874 297850 58350
rect 182 53702 297750 53874
rect 182 53034 297850 53702
rect 270 52862 297850 53034
rect 182 48274 297850 52862
rect 182 48102 297750 48274
rect 182 47546 297850 48102
rect 270 47374 297850 47546
rect 182 42674 297850 47374
rect 182 42502 297750 42674
rect 182 42058 297850 42502
rect 270 41886 297850 42058
rect 182 37074 297850 41886
rect 182 36902 297750 37074
rect 182 36570 297850 36902
rect 270 36398 297850 36570
rect 182 31474 297850 36398
rect 182 31302 297750 31474
rect 182 31082 297850 31302
rect 270 30910 297850 31082
rect 182 25874 297850 30910
rect 182 25702 297750 25874
rect 182 25594 297850 25702
rect 270 25422 297850 25594
rect 182 20274 297850 25422
rect 182 20106 297750 20274
rect 270 20102 297750 20106
rect 270 19934 297850 20102
rect 182 14674 297850 19934
rect 182 14618 297750 14674
rect 270 14502 297750 14618
rect 270 14446 297850 14502
rect 182 9130 297850 14446
rect 270 9074 297850 9130
rect 270 8958 297750 9074
rect 182 8902 297750 8958
rect 182 3642 297850 8902
rect 270 3474 297850 3642
rect 270 3470 297750 3474
rect 182 3302 297750 3470
rect 182 1918 297850 3302
<< metal4 >>
rect -958 -822 -648 299134
rect -478 -342 -168 298654
rect 1577 -822 1887 299134
rect 3437 -822 3747 299134
rect 10577 -822 10887 299134
rect 12437 -822 12747 299134
rect 19577 -822 19887 299134
rect 21437 -822 21747 299134
rect 28577 -822 28887 299134
rect 30437 -822 30747 299134
rect 37577 -822 37887 299134
rect 39437 -822 39747 299134
rect 46577 -822 46887 299134
rect 48437 -822 48747 299134
rect 55577 -822 55887 299134
rect 57437 -822 57747 299134
rect 64577 -822 64887 299134
rect 66437 -822 66747 299134
rect 73577 -822 73887 299134
rect 75437 -822 75747 299134
rect 82577 -822 82887 299134
rect 84437 -822 84747 299134
rect 91577 -822 91887 299134
rect 93437 -822 93747 299134
rect 100577 -822 100887 299134
rect 102437 -822 102747 299134
rect 109577 -822 109887 299134
rect 111437 -822 111747 299134
rect 118577 -822 118887 299134
rect 120437 -822 120747 299134
rect 127577 228466 127887 299134
rect 127577 -822 127887 169510
rect 129437 -822 129747 299134
rect 136577 -822 136887 299134
rect 138437 -822 138747 299134
rect 145577 228259 145887 299134
rect 147437 228259 147747 299134
rect 154577 228259 154887 299134
rect 156437 228259 156747 299134
rect 145577 -822 145887 223085
rect 147437 -822 147747 223085
rect 154577 -822 154887 223085
rect 156437 -822 156747 223085
rect 163577 -822 163887 299134
rect 165437 -822 165747 299134
rect 172577 -822 172887 299134
rect 174437 -822 174747 299134
rect 181577 -822 181887 299134
rect 183437 -822 183747 299134
rect 190577 -822 190887 299134
rect 192437 -822 192747 299134
rect 199577 -822 199887 299134
rect 201437 -822 201747 299134
rect 208577 -822 208887 299134
rect 210437 -822 210747 299134
rect 217577 -822 217887 299134
rect 219437 -822 219747 299134
rect 226577 -822 226887 299134
rect 228437 -822 228747 299134
rect 235577 -822 235887 299134
rect 237437 -822 237747 299134
rect 244577 -822 244887 299134
rect 246437 -822 246747 299134
rect 253577 -822 253887 299134
rect 255437 -822 255747 299134
rect 262577 -822 262887 299134
rect 264437 -822 264747 299134
rect 271577 -822 271887 299134
rect 273437 -822 273747 299134
rect 280577 -822 280887 299134
rect 282437 -822 282747 299134
rect 289577 -822 289887 299134
rect 291437 -822 291747 299134
rect 298200 -342 298510 298654
rect 298680 -822 298990 299134
<< obsm4 >>
rect 119724 170538 120407 228975
rect 120777 228436 127547 228975
rect 127917 228436 129407 228975
rect 120777 170538 129407 228436
rect 129777 170538 136547 228975
rect 136917 170538 138407 228975
rect 138777 228229 145547 228975
rect 145917 228229 147407 228975
rect 147777 228229 154547 228975
rect 154917 228229 156407 228975
rect 156777 228229 163547 228975
rect 138777 223115 163547 228229
rect 138777 170538 145547 223115
rect 145917 170538 147407 223115
rect 147777 170538 154547 223115
rect 154917 170538 156407 223115
rect 156777 170538 163547 223115
rect 163917 170538 165407 228975
rect 165777 170538 172547 228975
rect 172917 170538 173644 228975
<< metal5 >>
rect -958 298824 298990 299134
rect -478 298344 298510 298654
rect -958 292913 298990 293223
rect -958 289913 298990 290223
rect -958 283913 298990 284223
rect -958 280913 298990 281223
rect -958 274913 298990 275223
rect -958 271913 298990 272223
rect -958 265913 298990 266223
rect -958 262913 298990 263223
rect -958 256913 298990 257223
rect -958 253913 298990 254223
rect -958 247913 298990 248223
rect -958 244913 298990 245223
rect -958 238913 298990 239223
rect -958 235913 298990 236223
rect -958 229913 298990 230223
rect -958 226913 298990 227223
rect -958 220913 298990 221223
rect -958 217913 298990 218223
rect -958 211913 298990 212223
rect -958 208913 298990 209223
rect -958 202913 298990 203223
rect -958 199913 298990 200223
rect -958 193913 298990 194223
rect -958 190913 298990 191223
rect -958 184913 298990 185223
rect -958 181913 298990 182223
rect -958 175913 298990 176223
rect -958 172913 298990 173223
rect -958 166913 298990 167223
rect -958 163913 298990 164223
rect -958 157913 298990 158223
rect -958 154913 298990 155223
rect -958 148913 298990 149223
rect -958 145913 298990 146223
rect -958 139913 298990 140223
rect -958 136913 298990 137223
rect -958 130913 298990 131223
rect -958 127913 298990 128223
rect -958 121913 298990 122223
rect -958 118913 298990 119223
rect -958 112913 298990 113223
rect -958 109913 298990 110223
rect -958 103913 298990 104223
rect -958 100913 298990 101223
rect -958 94913 298990 95223
rect -958 91913 298990 92223
rect -958 85913 298990 86223
rect -958 82913 298990 83223
rect -958 76913 298990 77223
rect -958 73913 298990 74223
rect -958 67913 298990 68223
rect -958 64913 298990 65223
rect -958 58913 298990 59223
rect -958 55913 298990 56223
rect -958 49913 298990 50223
rect -958 46913 298990 47223
rect -958 40913 298990 41223
rect -958 37913 298990 38223
rect -958 31913 298990 32223
rect -958 28913 298990 29223
rect -958 22913 298990 23223
rect -958 19913 298990 20223
rect -958 13913 298990 14223
rect -958 10913 298990 11223
rect -958 4913 298990 5223
rect -958 1913 298990 2223
rect -478 -342 298510 -32
rect -958 -822 298990 -512
<< labels >>
rlabel metal3 s 297780 120932 298500 121044 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal2 s 227164 297780 227276 298500 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 194236 297780 194348 298500 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 161308 297780 161420 298500 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 128380 297780 128492 298500 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 95452 297780 95564 298500 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 62524 297780 62636 298500 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 29596 297780 29708 298500 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal3 s -480 294364 240 294476 4 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s -480 272412 240 272524 4 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal3 s -480 250460 240 250572 4 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 297780 143332 298500 143444 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s -480 228508 240 228620 4 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s -480 206556 240 206668 4 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s -480 184604 240 184716 4 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal3 s -480 162652 240 162764 4 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s -480 140700 240 140812 4 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s -480 118748 240 118860 4 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s -480 96796 240 96908 4 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s -480 74844 240 74956 4 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s -480 52892 240 53004 4 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 297780 165732 298500 165844 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 297780 188132 298500 188244 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal3 s 297780 210532 298500 210644 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 297780 232932 298500 233044 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal3 s 297780 255332 298500 255444 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal3 s 297780 277732 298500 277844 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 293020 297780 293132 298500 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal2 s 260092 297780 260204 298500 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal3 s 297780 3332 298500 3444 6 io_in[0]
port 30 nsew signal input
rlabel metal3 s 297780 193732 298500 193844 6 io_in[10]
port 31 nsew signal input
rlabel metal3 s 297780 216132 298500 216244 6 io_in[11]
port 32 nsew signal input
rlabel metal3 s 297780 238532 298500 238644 6 io_in[12]
port 33 nsew signal input
rlabel metal3 s 297780 260932 298500 261044 6 io_in[13]
port 34 nsew signal input
rlabel metal3 s 297780 283332 298500 283444 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 284788 297780 284900 298500 6 io_in[15]
port 36 nsew signal input
rlabel metal2 s 251860 297780 251972 298500 6 io_in[16]
port 37 nsew signal input
rlabel metal2 s 218932 297780 219044 298500 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 186004 297780 186116 298500 6 io_in[18]
port 39 nsew signal input
rlabel metal2 s 153076 297780 153188 298500 6 io_in[19]
port 40 nsew signal input
rlabel metal3 s 297780 20132 298500 20244 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 120148 297780 120260 298500 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 87220 297780 87332 298500 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 54292 297780 54404 298500 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 21364 297780 21476 298500 6 io_in[23]
port 45 nsew signal input
rlabel metal3 s -480 288876 240 288988 4 io_in[24]
port 46 nsew signal input
rlabel metal3 s -480 266924 240 267036 4 io_in[25]
port 47 nsew signal input
rlabel metal3 s -480 244972 240 245084 4 io_in[26]
port 48 nsew signal input
rlabel metal3 s -480 223020 240 223132 4 io_in[27]
port 49 nsew signal input
rlabel metal3 s -480 201068 240 201180 4 io_in[28]
port 50 nsew signal input
rlabel metal3 s -480 179116 240 179228 4 io_in[29]
port 51 nsew signal input
rlabel metal3 s 297780 36932 298500 37044 6 io_in[2]
port 52 nsew signal input
rlabel metal3 s -480 157164 240 157276 4 io_in[30]
port 53 nsew signal input
rlabel metal3 s -480 135212 240 135324 4 io_in[31]
port 54 nsew signal input
rlabel metal3 s -480 113260 240 113372 4 io_in[32]
port 55 nsew signal input
rlabel metal3 s -480 91308 240 91420 4 io_in[33]
port 56 nsew signal input
rlabel metal3 s -480 69356 240 69468 4 io_in[34]
port 57 nsew signal input
rlabel metal3 s -480 47404 240 47516 4 io_in[35]
port 58 nsew signal input
rlabel metal3 s -480 30940 240 31052 4 io_in[36]
port 59 nsew signal input
rlabel metal3 s -480 14476 240 14588 4 io_in[37]
port 60 nsew signal input
rlabel metal3 s 297780 53732 298500 53844 6 io_in[3]
port 61 nsew signal input
rlabel metal3 s 297780 70532 298500 70644 6 io_in[4]
port 62 nsew signal input
rlabel metal3 s 297780 87332 298500 87444 6 io_in[5]
port 63 nsew signal input
rlabel metal3 s 297780 104132 298500 104244 6 io_in[6]
port 64 nsew signal input
rlabel metal3 s 297780 126532 298500 126644 6 io_in[7]
port 65 nsew signal input
rlabel metal3 s 297780 148932 298500 149044 6 io_in[8]
port 66 nsew signal input
rlabel metal3 s 297780 171332 298500 171444 6 io_in[9]
port 67 nsew signal input
rlabel metal3 s 297780 14532 298500 14644 6 io_oeb[0]
port 68 nsew signal output
rlabel metal3 s 297780 204932 298500 205044 6 io_oeb[10]
port 69 nsew signal output
rlabel metal3 s 297780 227332 298500 227444 6 io_oeb[11]
port 70 nsew signal output
rlabel metal3 s 297780 249732 298500 249844 6 io_oeb[12]
port 71 nsew signal output
rlabel metal3 s 297780 272132 298500 272244 6 io_oeb[13]
port 72 nsew signal output
rlabel metal3 s 297780 294532 298500 294644 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 268324 297780 268436 298500 6 io_oeb[15]
port 74 nsew signal output
rlabel metal2 s 235396 297780 235508 298500 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 202468 297780 202580 298500 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 169540 297780 169652 298500 6 io_oeb[18]
port 77 nsew signal output
rlabel metal2 s 136612 297780 136724 298500 6 io_oeb[19]
port 78 nsew signal output
rlabel metal3 s 297780 31332 298500 31444 6 io_oeb[1]
port 79 nsew signal output
rlabel metal2 s 103684 297780 103796 298500 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 70756 297780 70868 298500 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 37828 297780 37940 298500 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 4900 297780 5012 298500 6 io_oeb[23]
port 83 nsew signal output
rlabel metal3 s -480 277900 240 278012 4 io_oeb[24]
port 84 nsew signal output
rlabel metal3 s -480 255948 240 256060 4 io_oeb[25]
port 85 nsew signal output
rlabel metal3 s -480 233996 240 234108 4 io_oeb[26]
port 86 nsew signal output
rlabel metal3 s -480 212044 240 212156 4 io_oeb[27]
port 87 nsew signal output
rlabel metal3 s -480 190092 240 190204 4 io_oeb[28]
port 88 nsew signal output
rlabel metal3 s -480 168140 240 168252 4 io_oeb[29]
port 89 nsew signal output
rlabel metal3 s 297780 48132 298500 48244 6 io_oeb[2]
port 90 nsew signal output
rlabel metal3 s -480 146188 240 146300 4 io_oeb[30]
port 91 nsew signal output
rlabel metal3 s -480 124236 240 124348 4 io_oeb[31]
port 92 nsew signal output
rlabel metal3 s -480 102284 240 102396 4 io_oeb[32]
port 93 nsew signal output
rlabel metal3 s -480 80332 240 80444 4 io_oeb[33]
port 94 nsew signal output
rlabel metal3 s -480 58380 240 58492 4 io_oeb[34]
port 95 nsew signal output
rlabel metal3 s -480 36428 240 36540 4 io_oeb[35]
port 96 nsew signal output
rlabel metal3 s -480 19964 240 20076 4 io_oeb[36]
port 97 nsew signal output
rlabel metal3 s -480 3500 240 3612 4 io_oeb[37]
port 98 nsew signal output
rlabel metal3 s 297780 64932 298500 65044 6 io_oeb[3]
port 99 nsew signal output
rlabel metal3 s 297780 81732 298500 81844 6 io_oeb[4]
port 100 nsew signal output
rlabel metal3 s 297780 98532 298500 98644 6 io_oeb[5]
port 101 nsew signal output
rlabel metal3 s 297780 115332 298500 115444 6 io_oeb[6]
port 102 nsew signal output
rlabel metal3 s 297780 137732 298500 137844 6 io_oeb[7]
port 103 nsew signal output
rlabel metal3 s 297780 160132 298500 160244 6 io_oeb[8]
port 104 nsew signal output
rlabel metal3 s 297780 182532 298500 182644 6 io_oeb[9]
port 105 nsew signal output
rlabel metal3 s 297780 8932 298500 9044 6 io_out[0]
port 106 nsew signal output
rlabel metal3 s 297780 199332 298500 199444 6 io_out[10]
port 107 nsew signal output
rlabel metal3 s 297780 221732 298500 221844 6 io_out[11]
port 108 nsew signal output
rlabel metal3 s 297780 244132 298500 244244 6 io_out[12]
port 109 nsew signal output
rlabel metal3 s 297780 266532 298500 266644 6 io_out[13]
port 110 nsew signal output
rlabel metal3 s 297780 288932 298500 289044 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 276556 297780 276668 298500 6 io_out[15]
port 112 nsew signal output
rlabel metal2 s 243628 297780 243740 298500 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 210700 297780 210812 298500 6 io_out[17]
port 114 nsew signal output
rlabel metal2 s 177772 297780 177884 298500 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 144844 297780 144956 298500 6 io_out[19]
port 116 nsew signal output
rlabel metal3 s 297780 25732 298500 25844 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 111916 297780 112028 298500 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 78988 297780 79100 298500 6 io_out[21]
port 119 nsew signal output
rlabel metal2 s 46060 297780 46172 298500 6 io_out[22]
port 120 nsew signal output
rlabel metal2 s 13132 297780 13244 298500 6 io_out[23]
port 121 nsew signal output
rlabel metal3 s -480 283388 240 283500 4 io_out[24]
port 122 nsew signal output
rlabel metal3 s -480 261436 240 261548 4 io_out[25]
port 123 nsew signal output
rlabel metal3 s -480 239484 240 239596 4 io_out[26]
port 124 nsew signal output
rlabel metal3 s -480 217532 240 217644 4 io_out[27]
port 125 nsew signal output
rlabel metal3 s -480 195580 240 195692 4 io_out[28]
port 126 nsew signal output
rlabel metal3 s -480 173628 240 173740 4 io_out[29]
port 127 nsew signal output
rlabel metal3 s 297780 42532 298500 42644 6 io_out[2]
port 128 nsew signal output
rlabel metal3 s -480 151676 240 151788 4 io_out[30]
port 129 nsew signal output
rlabel metal3 s -480 129724 240 129836 4 io_out[31]
port 130 nsew signal output
rlabel metal3 s -480 107772 240 107884 4 io_out[32]
port 131 nsew signal output
rlabel metal3 s -480 85820 240 85932 4 io_out[33]
port 132 nsew signal output
rlabel metal3 s -480 63868 240 63980 4 io_out[34]
port 133 nsew signal output
rlabel metal3 s -480 41916 240 42028 4 io_out[35]
port 134 nsew signal output
rlabel metal3 s -480 25452 240 25564 4 io_out[36]
port 135 nsew signal output
rlabel metal3 s -480 8988 240 9100 4 io_out[37]
port 136 nsew signal output
rlabel metal3 s 297780 59332 298500 59444 6 io_out[3]
port 137 nsew signal output
rlabel metal3 s 297780 76132 298500 76244 6 io_out[4]
port 138 nsew signal output
rlabel metal3 s 297780 92932 298500 93044 6 io_out[5]
port 139 nsew signal output
rlabel metal3 s 297780 109732 298500 109844 6 io_out[6]
port 140 nsew signal output
rlabel metal3 s 297780 132132 298500 132244 6 io_out[7]
port 141 nsew signal output
rlabel metal3 s 297780 154532 298500 154644 6 io_out[8]
port 142 nsew signal output
rlabel metal3 s 297780 176932 298500 177044 6 io_out[9]
port 143 nsew signal output
rlabel metal2 s 106596 -480 106708 240 8 la_data_in[0]
port 144 nsew signal input
rlabel metal2 s 135156 -480 135268 240 8 la_data_in[10]
port 145 nsew signal input
rlabel metal2 s 138012 -480 138124 240 8 la_data_in[11]
port 146 nsew signal input
rlabel metal2 s 140868 -480 140980 240 8 la_data_in[12]
port 147 nsew signal input
rlabel metal2 s 143724 -480 143836 240 8 la_data_in[13]
port 148 nsew signal input
rlabel metal2 s 146580 -480 146692 240 8 la_data_in[14]
port 149 nsew signal input
rlabel metal2 s 149436 -480 149548 240 8 la_data_in[15]
port 150 nsew signal input
rlabel metal2 s 152292 -480 152404 240 8 la_data_in[16]
port 151 nsew signal input
rlabel metal2 s 155148 -480 155260 240 8 la_data_in[17]
port 152 nsew signal input
rlabel metal2 s 158004 -480 158116 240 8 la_data_in[18]
port 153 nsew signal input
rlabel metal2 s 160860 -480 160972 240 8 la_data_in[19]
port 154 nsew signal input
rlabel metal2 s 109452 -480 109564 240 8 la_data_in[1]
port 155 nsew signal input
rlabel metal2 s 163716 -480 163828 240 8 la_data_in[20]
port 156 nsew signal input
rlabel metal2 s 166572 -480 166684 240 8 la_data_in[21]
port 157 nsew signal input
rlabel metal2 s 169428 -480 169540 240 8 la_data_in[22]
port 158 nsew signal input
rlabel metal2 s 172284 -480 172396 240 8 la_data_in[23]
port 159 nsew signal input
rlabel metal2 s 175140 -480 175252 240 8 la_data_in[24]
port 160 nsew signal input
rlabel metal2 s 177996 -480 178108 240 8 la_data_in[25]
port 161 nsew signal input
rlabel metal2 s 180852 -480 180964 240 8 la_data_in[26]
port 162 nsew signal input
rlabel metal2 s 183708 -480 183820 240 8 la_data_in[27]
port 163 nsew signal input
rlabel metal2 s 186564 -480 186676 240 8 la_data_in[28]
port 164 nsew signal input
rlabel metal2 s 189420 -480 189532 240 8 la_data_in[29]
port 165 nsew signal input
rlabel metal2 s 112308 -480 112420 240 8 la_data_in[2]
port 166 nsew signal input
rlabel metal2 s 192276 -480 192388 240 8 la_data_in[30]
port 167 nsew signal input
rlabel metal2 s 195132 -480 195244 240 8 la_data_in[31]
port 168 nsew signal input
rlabel metal2 s 197988 -480 198100 240 8 la_data_in[32]
port 169 nsew signal input
rlabel metal2 s 200844 -480 200956 240 8 la_data_in[33]
port 170 nsew signal input
rlabel metal2 s 203700 -480 203812 240 8 la_data_in[34]
port 171 nsew signal input
rlabel metal2 s 206556 -480 206668 240 8 la_data_in[35]
port 172 nsew signal input
rlabel metal2 s 209412 -480 209524 240 8 la_data_in[36]
port 173 nsew signal input
rlabel metal2 s 212268 -480 212380 240 8 la_data_in[37]
port 174 nsew signal input
rlabel metal2 s 215124 -480 215236 240 8 la_data_in[38]
port 175 nsew signal input
rlabel metal2 s 217980 -480 218092 240 8 la_data_in[39]
port 176 nsew signal input
rlabel metal2 s 115164 -480 115276 240 8 la_data_in[3]
port 177 nsew signal input
rlabel metal2 s 220836 -480 220948 240 8 la_data_in[40]
port 178 nsew signal input
rlabel metal2 s 223692 -480 223804 240 8 la_data_in[41]
port 179 nsew signal input
rlabel metal2 s 226548 -480 226660 240 8 la_data_in[42]
port 180 nsew signal input
rlabel metal2 s 229404 -480 229516 240 8 la_data_in[43]
port 181 nsew signal input
rlabel metal2 s 232260 -480 232372 240 8 la_data_in[44]
port 182 nsew signal input
rlabel metal2 s 235116 -480 235228 240 8 la_data_in[45]
port 183 nsew signal input
rlabel metal2 s 237972 -480 238084 240 8 la_data_in[46]
port 184 nsew signal input
rlabel metal2 s 240828 -480 240940 240 8 la_data_in[47]
port 185 nsew signal input
rlabel metal2 s 243684 -480 243796 240 8 la_data_in[48]
port 186 nsew signal input
rlabel metal2 s 246540 -480 246652 240 8 la_data_in[49]
port 187 nsew signal input
rlabel metal2 s 118020 -480 118132 240 8 la_data_in[4]
port 188 nsew signal input
rlabel metal2 s 249396 -480 249508 240 8 la_data_in[50]
port 189 nsew signal input
rlabel metal2 s 252252 -480 252364 240 8 la_data_in[51]
port 190 nsew signal input
rlabel metal2 s 255108 -480 255220 240 8 la_data_in[52]
port 191 nsew signal input
rlabel metal2 s 257964 -480 258076 240 8 la_data_in[53]
port 192 nsew signal input
rlabel metal2 s 260820 -480 260932 240 8 la_data_in[54]
port 193 nsew signal input
rlabel metal2 s 263676 -480 263788 240 8 la_data_in[55]
port 194 nsew signal input
rlabel metal2 s 266532 -480 266644 240 8 la_data_in[56]
port 195 nsew signal input
rlabel metal2 s 269388 -480 269500 240 8 la_data_in[57]
port 196 nsew signal input
rlabel metal2 s 272244 -480 272356 240 8 la_data_in[58]
port 197 nsew signal input
rlabel metal2 s 275100 -480 275212 240 8 la_data_in[59]
port 198 nsew signal input
rlabel metal2 s 120876 -480 120988 240 8 la_data_in[5]
port 199 nsew signal input
rlabel metal2 s 277956 -480 278068 240 8 la_data_in[60]
port 200 nsew signal input
rlabel metal2 s 280812 -480 280924 240 8 la_data_in[61]
port 201 nsew signal input
rlabel metal2 s 283668 -480 283780 240 8 la_data_in[62]
port 202 nsew signal input
rlabel metal2 s 286524 -480 286636 240 8 la_data_in[63]
port 203 nsew signal input
rlabel metal2 s 123732 -480 123844 240 8 la_data_in[6]
port 204 nsew signal input
rlabel metal2 s 126588 -480 126700 240 8 la_data_in[7]
port 205 nsew signal input
rlabel metal2 s 129444 -480 129556 240 8 la_data_in[8]
port 206 nsew signal input
rlabel metal2 s 132300 -480 132412 240 8 la_data_in[9]
port 207 nsew signal input
rlabel metal2 s 107548 -480 107660 240 8 la_data_out[0]
port 208 nsew signal output
rlabel metal2 s 136108 -480 136220 240 8 la_data_out[10]
port 209 nsew signal output
rlabel metal2 s 138964 -480 139076 240 8 la_data_out[11]
port 210 nsew signal output
rlabel metal2 s 141820 -480 141932 240 8 la_data_out[12]
port 211 nsew signal output
rlabel metal2 s 144676 -480 144788 240 8 la_data_out[13]
port 212 nsew signal output
rlabel metal2 s 147532 -480 147644 240 8 la_data_out[14]
port 213 nsew signal output
rlabel metal2 s 150388 -480 150500 240 8 la_data_out[15]
port 214 nsew signal output
rlabel metal2 s 153244 -480 153356 240 8 la_data_out[16]
port 215 nsew signal output
rlabel metal2 s 156100 -480 156212 240 8 la_data_out[17]
port 216 nsew signal output
rlabel metal2 s 158956 -480 159068 240 8 la_data_out[18]
port 217 nsew signal output
rlabel metal2 s 161812 -480 161924 240 8 la_data_out[19]
port 218 nsew signal output
rlabel metal2 s 110404 -480 110516 240 8 la_data_out[1]
port 219 nsew signal output
rlabel metal2 s 164668 -480 164780 240 8 la_data_out[20]
port 220 nsew signal output
rlabel metal2 s 167524 -480 167636 240 8 la_data_out[21]
port 221 nsew signal output
rlabel metal2 s 170380 -480 170492 240 8 la_data_out[22]
port 222 nsew signal output
rlabel metal2 s 173236 -480 173348 240 8 la_data_out[23]
port 223 nsew signal output
rlabel metal2 s 176092 -480 176204 240 8 la_data_out[24]
port 224 nsew signal output
rlabel metal2 s 178948 -480 179060 240 8 la_data_out[25]
port 225 nsew signal output
rlabel metal2 s 181804 -480 181916 240 8 la_data_out[26]
port 226 nsew signal output
rlabel metal2 s 184660 -480 184772 240 8 la_data_out[27]
port 227 nsew signal output
rlabel metal2 s 187516 -480 187628 240 8 la_data_out[28]
port 228 nsew signal output
rlabel metal2 s 190372 -480 190484 240 8 la_data_out[29]
port 229 nsew signal output
rlabel metal2 s 113260 -480 113372 240 8 la_data_out[2]
port 230 nsew signal output
rlabel metal2 s 193228 -480 193340 240 8 la_data_out[30]
port 231 nsew signal output
rlabel metal2 s 196084 -480 196196 240 8 la_data_out[31]
port 232 nsew signal output
rlabel metal2 s 198940 -480 199052 240 8 la_data_out[32]
port 233 nsew signal output
rlabel metal2 s 201796 -480 201908 240 8 la_data_out[33]
port 234 nsew signal output
rlabel metal2 s 204652 -480 204764 240 8 la_data_out[34]
port 235 nsew signal output
rlabel metal2 s 207508 -480 207620 240 8 la_data_out[35]
port 236 nsew signal output
rlabel metal2 s 210364 -480 210476 240 8 la_data_out[36]
port 237 nsew signal output
rlabel metal2 s 213220 -480 213332 240 8 la_data_out[37]
port 238 nsew signal output
rlabel metal2 s 216076 -480 216188 240 8 la_data_out[38]
port 239 nsew signal output
rlabel metal2 s 218932 -480 219044 240 8 la_data_out[39]
port 240 nsew signal output
rlabel metal2 s 116116 -480 116228 240 8 la_data_out[3]
port 241 nsew signal output
rlabel metal2 s 221788 -480 221900 240 8 la_data_out[40]
port 242 nsew signal output
rlabel metal2 s 224644 -480 224756 240 8 la_data_out[41]
port 243 nsew signal output
rlabel metal2 s 227500 -480 227612 240 8 la_data_out[42]
port 244 nsew signal output
rlabel metal2 s 230356 -480 230468 240 8 la_data_out[43]
port 245 nsew signal output
rlabel metal2 s 233212 -480 233324 240 8 la_data_out[44]
port 246 nsew signal output
rlabel metal2 s 236068 -480 236180 240 8 la_data_out[45]
port 247 nsew signal output
rlabel metal2 s 238924 -480 239036 240 8 la_data_out[46]
port 248 nsew signal output
rlabel metal2 s 241780 -480 241892 240 8 la_data_out[47]
port 249 nsew signal output
rlabel metal2 s 244636 -480 244748 240 8 la_data_out[48]
port 250 nsew signal output
rlabel metal2 s 247492 -480 247604 240 8 la_data_out[49]
port 251 nsew signal output
rlabel metal2 s 118972 -480 119084 240 8 la_data_out[4]
port 252 nsew signal output
rlabel metal2 s 250348 -480 250460 240 8 la_data_out[50]
port 253 nsew signal output
rlabel metal2 s 253204 -480 253316 240 8 la_data_out[51]
port 254 nsew signal output
rlabel metal2 s 256060 -480 256172 240 8 la_data_out[52]
port 255 nsew signal output
rlabel metal2 s 258916 -480 259028 240 8 la_data_out[53]
port 256 nsew signal output
rlabel metal2 s 261772 -480 261884 240 8 la_data_out[54]
port 257 nsew signal output
rlabel metal2 s 264628 -480 264740 240 8 la_data_out[55]
port 258 nsew signal output
rlabel metal2 s 267484 -480 267596 240 8 la_data_out[56]
port 259 nsew signal output
rlabel metal2 s 270340 -480 270452 240 8 la_data_out[57]
port 260 nsew signal output
rlabel metal2 s 273196 -480 273308 240 8 la_data_out[58]
port 261 nsew signal output
rlabel metal2 s 276052 -480 276164 240 8 la_data_out[59]
port 262 nsew signal output
rlabel metal2 s 121828 -480 121940 240 8 la_data_out[5]
port 263 nsew signal output
rlabel metal2 s 278908 -480 279020 240 8 la_data_out[60]
port 264 nsew signal output
rlabel metal2 s 281764 -480 281876 240 8 la_data_out[61]
port 265 nsew signal output
rlabel metal2 s 284620 -480 284732 240 8 la_data_out[62]
port 266 nsew signal output
rlabel metal2 s 287476 -480 287588 240 8 la_data_out[63]
port 267 nsew signal output
rlabel metal2 s 124684 -480 124796 240 8 la_data_out[6]
port 268 nsew signal output
rlabel metal2 s 127540 -480 127652 240 8 la_data_out[7]
port 269 nsew signal output
rlabel metal2 s 130396 -480 130508 240 8 la_data_out[8]
port 270 nsew signal output
rlabel metal2 s 133252 -480 133364 240 8 la_data_out[9]
port 271 nsew signal output
rlabel metal2 s 108500 -480 108612 240 8 la_oenb[0]
port 272 nsew signal input
rlabel metal2 s 137060 -480 137172 240 8 la_oenb[10]
port 273 nsew signal input
rlabel metal2 s 139916 -480 140028 240 8 la_oenb[11]
port 274 nsew signal input
rlabel metal2 s 142772 -480 142884 240 8 la_oenb[12]
port 275 nsew signal input
rlabel metal2 s 145628 -480 145740 240 8 la_oenb[13]
port 276 nsew signal input
rlabel metal2 s 148484 -480 148596 240 8 la_oenb[14]
port 277 nsew signal input
rlabel metal2 s 151340 -480 151452 240 8 la_oenb[15]
port 278 nsew signal input
rlabel metal2 s 154196 -480 154308 240 8 la_oenb[16]
port 279 nsew signal input
rlabel metal2 s 157052 -480 157164 240 8 la_oenb[17]
port 280 nsew signal input
rlabel metal2 s 159908 -480 160020 240 8 la_oenb[18]
port 281 nsew signal input
rlabel metal2 s 162764 -480 162876 240 8 la_oenb[19]
port 282 nsew signal input
rlabel metal2 s 111356 -480 111468 240 8 la_oenb[1]
port 283 nsew signal input
rlabel metal2 s 165620 -480 165732 240 8 la_oenb[20]
port 284 nsew signal input
rlabel metal2 s 168476 -480 168588 240 8 la_oenb[21]
port 285 nsew signal input
rlabel metal2 s 171332 -480 171444 240 8 la_oenb[22]
port 286 nsew signal input
rlabel metal2 s 174188 -480 174300 240 8 la_oenb[23]
port 287 nsew signal input
rlabel metal2 s 177044 -480 177156 240 8 la_oenb[24]
port 288 nsew signal input
rlabel metal2 s 179900 -480 180012 240 8 la_oenb[25]
port 289 nsew signal input
rlabel metal2 s 182756 -480 182868 240 8 la_oenb[26]
port 290 nsew signal input
rlabel metal2 s 185612 -480 185724 240 8 la_oenb[27]
port 291 nsew signal input
rlabel metal2 s 188468 -480 188580 240 8 la_oenb[28]
port 292 nsew signal input
rlabel metal2 s 191324 -480 191436 240 8 la_oenb[29]
port 293 nsew signal input
rlabel metal2 s 114212 -480 114324 240 8 la_oenb[2]
port 294 nsew signal input
rlabel metal2 s 194180 -480 194292 240 8 la_oenb[30]
port 295 nsew signal input
rlabel metal2 s 197036 -480 197148 240 8 la_oenb[31]
port 296 nsew signal input
rlabel metal2 s 199892 -480 200004 240 8 la_oenb[32]
port 297 nsew signal input
rlabel metal2 s 202748 -480 202860 240 8 la_oenb[33]
port 298 nsew signal input
rlabel metal2 s 205604 -480 205716 240 8 la_oenb[34]
port 299 nsew signal input
rlabel metal2 s 208460 -480 208572 240 8 la_oenb[35]
port 300 nsew signal input
rlabel metal2 s 211316 -480 211428 240 8 la_oenb[36]
port 301 nsew signal input
rlabel metal2 s 214172 -480 214284 240 8 la_oenb[37]
port 302 nsew signal input
rlabel metal2 s 217028 -480 217140 240 8 la_oenb[38]
port 303 nsew signal input
rlabel metal2 s 219884 -480 219996 240 8 la_oenb[39]
port 304 nsew signal input
rlabel metal2 s 117068 -480 117180 240 8 la_oenb[3]
port 305 nsew signal input
rlabel metal2 s 222740 -480 222852 240 8 la_oenb[40]
port 306 nsew signal input
rlabel metal2 s 225596 -480 225708 240 8 la_oenb[41]
port 307 nsew signal input
rlabel metal2 s 228452 -480 228564 240 8 la_oenb[42]
port 308 nsew signal input
rlabel metal2 s 231308 -480 231420 240 8 la_oenb[43]
port 309 nsew signal input
rlabel metal2 s 234164 -480 234276 240 8 la_oenb[44]
port 310 nsew signal input
rlabel metal2 s 237020 -480 237132 240 8 la_oenb[45]
port 311 nsew signal input
rlabel metal2 s 239876 -480 239988 240 8 la_oenb[46]
port 312 nsew signal input
rlabel metal2 s 242732 -480 242844 240 8 la_oenb[47]
port 313 nsew signal input
rlabel metal2 s 245588 -480 245700 240 8 la_oenb[48]
port 314 nsew signal input
rlabel metal2 s 248444 -480 248556 240 8 la_oenb[49]
port 315 nsew signal input
rlabel metal2 s 119924 -480 120036 240 8 la_oenb[4]
port 316 nsew signal input
rlabel metal2 s 251300 -480 251412 240 8 la_oenb[50]
port 317 nsew signal input
rlabel metal2 s 254156 -480 254268 240 8 la_oenb[51]
port 318 nsew signal input
rlabel metal2 s 257012 -480 257124 240 8 la_oenb[52]
port 319 nsew signal input
rlabel metal2 s 259868 -480 259980 240 8 la_oenb[53]
port 320 nsew signal input
rlabel metal2 s 262724 -480 262836 240 8 la_oenb[54]
port 321 nsew signal input
rlabel metal2 s 265580 -480 265692 240 8 la_oenb[55]
port 322 nsew signal input
rlabel metal2 s 268436 -480 268548 240 8 la_oenb[56]
port 323 nsew signal input
rlabel metal2 s 271292 -480 271404 240 8 la_oenb[57]
port 324 nsew signal input
rlabel metal2 s 274148 -480 274260 240 8 la_oenb[58]
port 325 nsew signal input
rlabel metal2 s 277004 -480 277116 240 8 la_oenb[59]
port 326 nsew signal input
rlabel metal2 s 122780 -480 122892 240 8 la_oenb[5]
port 327 nsew signal input
rlabel metal2 s 279860 -480 279972 240 8 la_oenb[60]
port 328 nsew signal input
rlabel metal2 s 282716 -480 282828 240 8 la_oenb[61]
port 329 nsew signal input
rlabel metal2 s 285572 -480 285684 240 8 la_oenb[62]
port 330 nsew signal input
rlabel metal2 s 288428 -480 288540 240 8 la_oenb[63]
port 331 nsew signal input
rlabel metal2 s 125636 -480 125748 240 8 la_oenb[6]
port 332 nsew signal input
rlabel metal2 s 128492 -480 128604 240 8 la_oenb[7]
port 333 nsew signal input
rlabel metal2 s 131348 -480 131460 240 8 la_oenb[8]
port 334 nsew signal input
rlabel metal2 s 134204 -480 134316 240 8 la_oenb[9]
port 335 nsew signal input
rlabel metal2 s 289380 -480 289492 240 8 user_clock2
port 336 nsew signal input
rlabel metal2 s 290332 -480 290444 240 8 user_irq[0]
port 337 nsew signal output
rlabel metal2 s 291284 -480 291396 240 8 user_irq[1]
port 338 nsew signal output
rlabel metal2 s 292236 -480 292348 240 8 user_irq[2]
port 339 nsew signal output
rlabel metal4 s -478 -342 -168 298654 4 vdd
port 340 nsew power bidirectional
rlabel metal5 s -478 -342 298510 -32 8 vdd
port 340 nsew power bidirectional
rlabel metal5 s -478 298344 298510 298654 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 298200 -342 298510 298654 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 1577 -822 1887 299134 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 10577 -822 10887 299134 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 19577 -822 19887 299134 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 28577 -822 28887 299134 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 37577 -822 37887 299134 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 46577 -822 46887 299134 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 55577 -822 55887 299134 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 64577 -822 64887 299134 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 73577 -822 73887 299134 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 82577 -822 82887 299134 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 91577 -822 91887 299134 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 100577 -822 100887 299134 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 109577 -822 109887 299134 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 118577 -822 118887 299134 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 127577 -822 127887 169510 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 127577 228466 127887 299134 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 136577 -822 136887 299134 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 145577 -822 145887 223085 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 145577 228259 145887 299134 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 154577 -822 154887 223085 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 154577 228259 154887 299134 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 163577 -822 163887 299134 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 172577 -822 172887 299134 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 181577 -822 181887 299134 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 190577 -822 190887 299134 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 199577 -822 199887 299134 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 208577 -822 208887 299134 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 217577 -822 217887 299134 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 226577 -822 226887 299134 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 235577 -822 235887 299134 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 244577 -822 244887 299134 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 253577 -822 253887 299134 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 262577 -822 262887 299134 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 271577 -822 271887 299134 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 280577 -822 280887 299134 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 289577 -822 289887 299134 6 vdd
port 340 nsew power bidirectional
rlabel metal5 s -958 1913 298990 2223 6 vdd
port 340 nsew power bidirectional
rlabel metal5 s -958 10913 298990 11223 6 vdd
port 340 nsew power bidirectional
rlabel metal5 s -958 19913 298990 20223 6 vdd
port 340 nsew power bidirectional
rlabel metal5 s -958 28913 298990 29223 6 vdd
port 340 nsew power bidirectional
rlabel metal5 s -958 37913 298990 38223 6 vdd
port 340 nsew power bidirectional
rlabel metal5 s -958 46913 298990 47223 6 vdd
port 340 nsew power bidirectional
rlabel metal5 s -958 55913 298990 56223 6 vdd
port 340 nsew power bidirectional
rlabel metal5 s -958 64913 298990 65223 6 vdd
port 340 nsew power bidirectional
rlabel metal5 s -958 73913 298990 74223 6 vdd
port 340 nsew power bidirectional
rlabel metal5 s -958 82913 298990 83223 6 vdd
port 340 nsew power bidirectional
rlabel metal5 s -958 91913 298990 92223 6 vdd
port 340 nsew power bidirectional
rlabel metal5 s -958 100913 298990 101223 6 vdd
port 340 nsew power bidirectional
rlabel metal5 s -958 109913 298990 110223 6 vdd
port 340 nsew power bidirectional
rlabel metal5 s -958 118913 298990 119223 6 vdd
port 340 nsew power bidirectional
rlabel metal5 s -958 127913 298990 128223 6 vdd
port 340 nsew power bidirectional
rlabel metal5 s -958 136913 298990 137223 6 vdd
port 340 nsew power bidirectional
rlabel metal5 s -958 145913 298990 146223 6 vdd
port 340 nsew power bidirectional
rlabel metal5 s -958 154913 298990 155223 6 vdd
port 340 nsew power bidirectional
rlabel metal5 s -958 163913 298990 164223 6 vdd
port 340 nsew power bidirectional
rlabel metal5 s -958 172913 298990 173223 6 vdd
port 340 nsew power bidirectional
rlabel metal5 s -958 181913 298990 182223 6 vdd
port 340 nsew power bidirectional
rlabel metal5 s -958 190913 298990 191223 6 vdd
port 340 nsew power bidirectional
rlabel metal5 s -958 199913 298990 200223 6 vdd
port 340 nsew power bidirectional
rlabel metal5 s -958 208913 298990 209223 6 vdd
port 340 nsew power bidirectional
rlabel metal5 s -958 217913 298990 218223 6 vdd
port 340 nsew power bidirectional
rlabel metal5 s -958 226913 298990 227223 6 vdd
port 340 nsew power bidirectional
rlabel metal5 s -958 235913 298990 236223 6 vdd
port 340 nsew power bidirectional
rlabel metal5 s -958 244913 298990 245223 6 vdd
port 340 nsew power bidirectional
rlabel metal5 s -958 253913 298990 254223 6 vdd
port 340 nsew power bidirectional
rlabel metal5 s -958 262913 298990 263223 6 vdd
port 340 nsew power bidirectional
rlabel metal5 s -958 271913 298990 272223 6 vdd
port 340 nsew power bidirectional
rlabel metal5 s -958 280913 298990 281223 6 vdd
port 340 nsew power bidirectional
rlabel metal5 s -958 289913 298990 290223 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s -958 -822 -648 299134 4 vss
port 341 nsew ground bidirectional
rlabel metal5 s -958 -822 298990 -512 8 vss
port 341 nsew ground bidirectional
rlabel metal5 s -958 298824 298990 299134 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 298680 -822 298990 299134 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 3437 -822 3747 299134 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 12437 -822 12747 299134 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 21437 -822 21747 299134 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 30437 -822 30747 299134 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 39437 -822 39747 299134 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 48437 -822 48747 299134 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 57437 -822 57747 299134 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 66437 -822 66747 299134 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 75437 -822 75747 299134 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 84437 -822 84747 299134 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 93437 -822 93747 299134 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 102437 -822 102747 299134 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 111437 -822 111747 299134 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 120437 -822 120747 299134 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 129437 -822 129747 299134 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 138437 -822 138747 299134 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 147437 -822 147747 223085 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 147437 228259 147747 299134 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 156437 -822 156747 223085 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 156437 228259 156747 299134 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 165437 -822 165747 299134 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 174437 -822 174747 299134 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 183437 -822 183747 299134 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 192437 -822 192747 299134 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 201437 -822 201747 299134 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 210437 -822 210747 299134 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 219437 -822 219747 299134 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 228437 -822 228747 299134 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 237437 -822 237747 299134 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 246437 -822 246747 299134 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 255437 -822 255747 299134 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 264437 -822 264747 299134 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 273437 -822 273747 299134 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 282437 -822 282747 299134 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 291437 -822 291747 299134 6 vss
port 341 nsew ground bidirectional
rlabel metal5 s -958 4913 298990 5223 6 vss
port 341 nsew ground bidirectional
rlabel metal5 s -958 13913 298990 14223 6 vss
port 341 nsew ground bidirectional
rlabel metal5 s -958 22913 298990 23223 6 vss
port 341 nsew ground bidirectional
rlabel metal5 s -958 31913 298990 32223 6 vss
port 341 nsew ground bidirectional
rlabel metal5 s -958 40913 298990 41223 6 vss
port 341 nsew ground bidirectional
rlabel metal5 s -958 49913 298990 50223 6 vss
port 341 nsew ground bidirectional
rlabel metal5 s -958 58913 298990 59223 6 vss
port 341 nsew ground bidirectional
rlabel metal5 s -958 67913 298990 68223 6 vss
port 341 nsew ground bidirectional
rlabel metal5 s -958 76913 298990 77223 6 vss
port 341 nsew ground bidirectional
rlabel metal5 s -958 85913 298990 86223 6 vss
port 341 nsew ground bidirectional
rlabel metal5 s -958 94913 298990 95223 6 vss
port 341 nsew ground bidirectional
rlabel metal5 s -958 103913 298990 104223 6 vss
port 341 nsew ground bidirectional
rlabel metal5 s -958 112913 298990 113223 6 vss
port 341 nsew ground bidirectional
rlabel metal5 s -958 121913 298990 122223 6 vss
port 341 nsew ground bidirectional
rlabel metal5 s -958 130913 298990 131223 6 vss
port 341 nsew ground bidirectional
rlabel metal5 s -958 139913 298990 140223 6 vss
port 341 nsew ground bidirectional
rlabel metal5 s -958 148913 298990 149223 6 vss
port 341 nsew ground bidirectional
rlabel metal5 s -958 157913 298990 158223 6 vss
port 341 nsew ground bidirectional
rlabel metal5 s -958 166913 298990 167223 6 vss
port 341 nsew ground bidirectional
rlabel metal5 s -958 175913 298990 176223 6 vss
port 341 nsew ground bidirectional
rlabel metal5 s -958 184913 298990 185223 6 vss
port 341 nsew ground bidirectional
rlabel metal5 s -958 193913 298990 194223 6 vss
port 341 nsew ground bidirectional
rlabel metal5 s -958 202913 298990 203223 6 vss
port 341 nsew ground bidirectional
rlabel metal5 s -958 211913 298990 212223 6 vss
port 341 nsew ground bidirectional
rlabel metal5 s -958 220913 298990 221223 6 vss
port 341 nsew ground bidirectional
rlabel metal5 s -958 229913 298990 230223 6 vss
port 341 nsew ground bidirectional
rlabel metal5 s -958 238913 298990 239223 6 vss
port 341 nsew ground bidirectional
rlabel metal5 s -958 247913 298990 248223 6 vss
port 341 nsew ground bidirectional
rlabel metal5 s -958 256913 298990 257223 6 vss
port 341 nsew ground bidirectional
rlabel metal5 s -958 265913 298990 266223 6 vss
port 341 nsew ground bidirectional
rlabel metal5 s -958 274913 298990 275223 6 vss
port 341 nsew ground bidirectional
rlabel metal5 s -958 283913 298990 284223 6 vss
port 341 nsew ground bidirectional
rlabel metal5 s -958 292913 298990 293223 6 vss
port 341 nsew ground bidirectional
rlabel metal2 s 5684 -480 5796 240 8 wb_clk_i
port 342 nsew signal input
rlabel metal2 s 6636 -480 6748 240 8 wb_rst_i
port 343 nsew signal input
rlabel metal2 s 7588 -480 7700 240 8 wbs_ack_o
port 344 nsew signal output
rlabel metal2 s 11396 -480 11508 240 8 wbs_adr_i[0]
port 345 nsew signal input
rlabel metal2 s 43764 -480 43876 240 8 wbs_adr_i[10]
port 346 nsew signal input
rlabel metal2 s 46620 -480 46732 240 8 wbs_adr_i[11]
port 347 nsew signal input
rlabel metal2 s 49476 -480 49588 240 8 wbs_adr_i[12]
port 348 nsew signal input
rlabel metal2 s 52332 -480 52444 240 8 wbs_adr_i[13]
port 349 nsew signal input
rlabel metal2 s 55188 -480 55300 240 8 wbs_adr_i[14]
port 350 nsew signal input
rlabel metal2 s 58044 -480 58156 240 8 wbs_adr_i[15]
port 351 nsew signal input
rlabel metal2 s 60900 -480 61012 240 8 wbs_adr_i[16]
port 352 nsew signal input
rlabel metal2 s 63756 -480 63868 240 8 wbs_adr_i[17]
port 353 nsew signal input
rlabel metal2 s 66612 -480 66724 240 8 wbs_adr_i[18]
port 354 nsew signal input
rlabel metal2 s 69468 -480 69580 240 8 wbs_adr_i[19]
port 355 nsew signal input
rlabel metal2 s 15204 -480 15316 240 8 wbs_adr_i[1]
port 356 nsew signal input
rlabel metal2 s 72324 -480 72436 240 8 wbs_adr_i[20]
port 357 nsew signal input
rlabel metal2 s 75180 -480 75292 240 8 wbs_adr_i[21]
port 358 nsew signal input
rlabel metal2 s 78036 -480 78148 240 8 wbs_adr_i[22]
port 359 nsew signal input
rlabel metal2 s 80892 -480 81004 240 8 wbs_adr_i[23]
port 360 nsew signal input
rlabel metal2 s 83748 -480 83860 240 8 wbs_adr_i[24]
port 361 nsew signal input
rlabel metal2 s 86604 -480 86716 240 8 wbs_adr_i[25]
port 362 nsew signal input
rlabel metal2 s 89460 -480 89572 240 8 wbs_adr_i[26]
port 363 nsew signal input
rlabel metal2 s 92316 -480 92428 240 8 wbs_adr_i[27]
port 364 nsew signal input
rlabel metal2 s 95172 -480 95284 240 8 wbs_adr_i[28]
port 365 nsew signal input
rlabel metal2 s 98028 -480 98140 240 8 wbs_adr_i[29]
port 366 nsew signal input
rlabel metal2 s 19012 -480 19124 240 8 wbs_adr_i[2]
port 367 nsew signal input
rlabel metal2 s 100884 -480 100996 240 8 wbs_adr_i[30]
port 368 nsew signal input
rlabel metal2 s 103740 -480 103852 240 8 wbs_adr_i[31]
port 369 nsew signal input
rlabel metal2 s 22820 -480 22932 240 8 wbs_adr_i[3]
port 370 nsew signal input
rlabel metal2 s 26628 -480 26740 240 8 wbs_adr_i[4]
port 371 nsew signal input
rlabel metal2 s 29484 -480 29596 240 8 wbs_adr_i[5]
port 372 nsew signal input
rlabel metal2 s 32340 -480 32452 240 8 wbs_adr_i[6]
port 373 nsew signal input
rlabel metal2 s 35196 -480 35308 240 8 wbs_adr_i[7]
port 374 nsew signal input
rlabel metal2 s 38052 -480 38164 240 8 wbs_adr_i[8]
port 375 nsew signal input
rlabel metal2 s 40908 -480 41020 240 8 wbs_adr_i[9]
port 376 nsew signal input
rlabel metal2 s 8540 -480 8652 240 8 wbs_cyc_i
port 377 nsew signal input
rlabel metal2 s 12348 -480 12460 240 8 wbs_dat_i[0]
port 378 nsew signal input
rlabel metal2 s 44716 -480 44828 240 8 wbs_dat_i[10]
port 379 nsew signal input
rlabel metal2 s 47572 -480 47684 240 8 wbs_dat_i[11]
port 380 nsew signal input
rlabel metal2 s 50428 -480 50540 240 8 wbs_dat_i[12]
port 381 nsew signal input
rlabel metal2 s 53284 -480 53396 240 8 wbs_dat_i[13]
port 382 nsew signal input
rlabel metal2 s 56140 -480 56252 240 8 wbs_dat_i[14]
port 383 nsew signal input
rlabel metal2 s 58996 -480 59108 240 8 wbs_dat_i[15]
port 384 nsew signal input
rlabel metal2 s 61852 -480 61964 240 8 wbs_dat_i[16]
port 385 nsew signal input
rlabel metal2 s 64708 -480 64820 240 8 wbs_dat_i[17]
port 386 nsew signal input
rlabel metal2 s 67564 -480 67676 240 8 wbs_dat_i[18]
port 387 nsew signal input
rlabel metal2 s 70420 -480 70532 240 8 wbs_dat_i[19]
port 388 nsew signal input
rlabel metal2 s 16156 -480 16268 240 8 wbs_dat_i[1]
port 389 nsew signal input
rlabel metal2 s 73276 -480 73388 240 8 wbs_dat_i[20]
port 390 nsew signal input
rlabel metal2 s 76132 -480 76244 240 8 wbs_dat_i[21]
port 391 nsew signal input
rlabel metal2 s 78988 -480 79100 240 8 wbs_dat_i[22]
port 392 nsew signal input
rlabel metal2 s 81844 -480 81956 240 8 wbs_dat_i[23]
port 393 nsew signal input
rlabel metal2 s 84700 -480 84812 240 8 wbs_dat_i[24]
port 394 nsew signal input
rlabel metal2 s 87556 -480 87668 240 8 wbs_dat_i[25]
port 395 nsew signal input
rlabel metal2 s 90412 -480 90524 240 8 wbs_dat_i[26]
port 396 nsew signal input
rlabel metal2 s 93268 -480 93380 240 8 wbs_dat_i[27]
port 397 nsew signal input
rlabel metal2 s 96124 -480 96236 240 8 wbs_dat_i[28]
port 398 nsew signal input
rlabel metal2 s 98980 -480 99092 240 8 wbs_dat_i[29]
port 399 nsew signal input
rlabel metal2 s 19964 -480 20076 240 8 wbs_dat_i[2]
port 400 nsew signal input
rlabel metal2 s 101836 -480 101948 240 8 wbs_dat_i[30]
port 401 nsew signal input
rlabel metal2 s 104692 -480 104804 240 8 wbs_dat_i[31]
port 402 nsew signal input
rlabel metal2 s 23772 -480 23884 240 8 wbs_dat_i[3]
port 403 nsew signal input
rlabel metal2 s 27580 -480 27692 240 8 wbs_dat_i[4]
port 404 nsew signal input
rlabel metal2 s 30436 -480 30548 240 8 wbs_dat_i[5]
port 405 nsew signal input
rlabel metal2 s 33292 -480 33404 240 8 wbs_dat_i[6]
port 406 nsew signal input
rlabel metal2 s 36148 -480 36260 240 8 wbs_dat_i[7]
port 407 nsew signal input
rlabel metal2 s 39004 -480 39116 240 8 wbs_dat_i[8]
port 408 nsew signal input
rlabel metal2 s 41860 -480 41972 240 8 wbs_dat_i[9]
port 409 nsew signal input
rlabel metal2 s 13300 -480 13412 240 8 wbs_dat_o[0]
port 410 nsew signal output
rlabel metal2 s 45668 -480 45780 240 8 wbs_dat_o[10]
port 411 nsew signal output
rlabel metal2 s 48524 -480 48636 240 8 wbs_dat_o[11]
port 412 nsew signal output
rlabel metal2 s 51380 -480 51492 240 8 wbs_dat_o[12]
port 413 nsew signal output
rlabel metal2 s 54236 -480 54348 240 8 wbs_dat_o[13]
port 414 nsew signal output
rlabel metal2 s 57092 -480 57204 240 8 wbs_dat_o[14]
port 415 nsew signal output
rlabel metal2 s 59948 -480 60060 240 8 wbs_dat_o[15]
port 416 nsew signal output
rlabel metal2 s 62804 -480 62916 240 8 wbs_dat_o[16]
port 417 nsew signal output
rlabel metal2 s 65660 -480 65772 240 8 wbs_dat_o[17]
port 418 nsew signal output
rlabel metal2 s 68516 -480 68628 240 8 wbs_dat_o[18]
port 419 nsew signal output
rlabel metal2 s 71372 -480 71484 240 8 wbs_dat_o[19]
port 420 nsew signal output
rlabel metal2 s 17108 -480 17220 240 8 wbs_dat_o[1]
port 421 nsew signal output
rlabel metal2 s 74228 -480 74340 240 8 wbs_dat_o[20]
port 422 nsew signal output
rlabel metal2 s 77084 -480 77196 240 8 wbs_dat_o[21]
port 423 nsew signal output
rlabel metal2 s 79940 -480 80052 240 8 wbs_dat_o[22]
port 424 nsew signal output
rlabel metal2 s 82796 -480 82908 240 8 wbs_dat_o[23]
port 425 nsew signal output
rlabel metal2 s 85652 -480 85764 240 8 wbs_dat_o[24]
port 426 nsew signal output
rlabel metal2 s 88508 -480 88620 240 8 wbs_dat_o[25]
port 427 nsew signal output
rlabel metal2 s 91364 -480 91476 240 8 wbs_dat_o[26]
port 428 nsew signal output
rlabel metal2 s 94220 -480 94332 240 8 wbs_dat_o[27]
port 429 nsew signal output
rlabel metal2 s 97076 -480 97188 240 8 wbs_dat_o[28]
port 430 nsew signal output
rlabel metal2 s 99932 -480 100044 240 8 wbs_dat_o[29]
port 431 nsew signal output
rlabel metal2 s 20916 -480 21028 240 8 wbs_dat_o[2]
port 432 nsew signal output
rlabel metal2 s 102788 -480 102900 240 8 wbs_dat_o[30]
port 433 nsew signal output
rlabel metal2 s 105644 -480 105756 240 8 wbs_dat_o[31]
port 434 nsew signal output
rlabel metal2 s 24724 -480 24836 240 8 wbs_dat_o[3]
port 435 nsew signal output
rlabel metal2 s 28532 -480 28644 240 8 wbs_dat_o[4]
port 436 nsew signal output
rlabel metal2 s 31388 -480 31500 240 8 wbs_dat_o[5]
port 437 nsew signal output
rlabel metal2 s 34244 -480 34356 240 8 wbs_dat_o[6]
port 438 nsew signal output
rlabel metal2 s 37100 -480 37212 240 8 wbs_dat_o[7]
port 439 nsew signal output
rlabel metal2 s 39956 -480 40068 240 8 wbs_dat_o[8]
port 440 nsew signal output
rlabel metal2 s 42812 -480 42924 240 8 wbs_dat_o[9]
port 441 nsew signal output
rlabel metal2 s 14252 -480 14364 240 8 wbs_sel_i[0]
port 442 nsew signal input
rlabel metal2 s 18060 -480 18172 240 8 wbs_sel_i[1]
port 443 nsew signal input
rlabel metal2 s 21868 -480 21980 240 8 wbs_sel_i[2]
port 444 nsew signal input
rlabel metal2 s 25676 -480 25788 240 8 wbs_sel_i[3]
port 445 nsew signal input
rlabel metal2 s 9492 -480 9604 240 8 wbs_stb_i
port 446 nsew signal input
rlabel metal2 s 10444 -480 10556 240 8 wbs_we_i
port 447 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 298020 298020
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 4801904
string GDS_FILE /opt/caravel_180/openlane/user_project_wrapper/runs/22_12_05_07_28/results/signoff/user_project_wrapper.magic.gds
string GDS_START 1836024
<< end >>

