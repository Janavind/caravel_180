magic
tech gf180mcuC
magscale 1 5
timestamp 1670241674
<< obsm1 >>
rect 672 855 59304 58673
<< metal2 >>
rect 1232 59600 1288 60000
rect 1736 59600 1792 60000
rect 2240 59600 2296 60000
rect 2744 59600 2800 60000
rect 3248 59600 3304 60000
rect 3752 59600 3808 60000
rect 4256 59600 4312 60000
rect 4760 59600 4816 60000
rect 5264 59600 5320 60000
rect 5768 59600 5824 60000
rect 6272 59600 6328 60000
rect 6776 59600 6832 60000
rect 7280 59600 7336 60000
rect 7784 59600 7840 60000
rect 8288 59600 8344 60000
rect 8792 59600 8848 60000
rect 9296 59600 9352 60000
rect 9800 59600 9856 60000
rect 10304 59600 10360 60000
rect 10808 59600 10864 60000
rect 11312 59600 11368 60000
rect 11816 59600 11872 60000
rect 12320 59600 12376 60000
rect 12824 59600 12880 60000
rect 13328 59600 13384 60000
rect 13832 59600 13888 60000
rect 14336 59600 14392 60000
rect 14840 59600 14896 60000
rect 15344 59600 15400 60000
rect 15848 59600 15904 60000
rect 16352 59600 16408 60000
rect 16856 59600 16912 60000
rect 17360 59600 17416 60000
rect 17864 59600 17920 60000
rect 18368 59600 18424 60000
rect 18872 59600 18928 60000
rect 19376 59600 19432 60000
rect 19880 59600 19936 60000
rect 20384 59600 20440 60000
rect 20888 59600 20944 60000
rect 21392 59600 21448 60000
rect 21896 59600 21952 60000
rect 22400 59600 22456 60000
rect 22904 59600 22960 60000
rect 23408 59600 23464 60000
rect 23912 59600 23968 60000
rect 24416 59600 24472 60000
rect 24920 59600 24976 60000
rect 25424 59600 25480 60000
rect 25928 59600 25984 60000
rect 26432 59600 26488 60000
rect 26936 59600 26992 60000
rect 27440 59600 27496 60000
rect 27944 59600 28000 60000
rect 28448 59600 28504 60000
rect 28952 59600 29008 60000
rect 29456 59600 29512 60000
rect 29960 59600 30016 60000
rect 30464 59600 30520 60000
rect 30968 59600 31024 60000
rect 31472 59600 31528 60000
rect 31976 59600 32032 60000
rect 32480 59600 32536 60000
rect 32984 59600 33040 60000
rect 33488 59600 33544 60000
rect 33992 59600 34048 60000
rect 34496 59600 34552 60000
rect 35000 59600 35056 60000
rect 35504 59600 35560 60000
rect 36008 59600 36064 60000
rect 36512 59600 36568 60000
rect 37016 59600 37072 60000
rect 37520 59600 37576 60000
rect 38024 59600 38080 60000
rect 38528 59600 38584 60000
rect 39032 59600 39088 60000
rect 39536 59600 39592 60000
rect 40040 59600 40096 60000
rect 40544 59600 40600 60000
rect 41048 59600 41104 60000
rect 41552 59600 41608 60000
rect 42056 59600 42112 60000
rect 42560 59600 42616 60000
rect 43064 59600 43120 60000
rect 43568 59600 43624 60000
rect 44072 59600 44128 60000
rect 44576 59600 44632 60000
rect 45080 59600 45136 60000
rect 45584 59600 45640 60000
rect 46088 59600 46144 60000
rect 46592 59600 46648 60000
rect 47096 59600 47152 60000
rect 47600 59600 47656 60000
rect 48104 59600 48160 60000
rect 48608 59600 48664 60000
rect 49112 59600 49168 60000
rect 49616 59600 49672 60000
rect 50120 59600 50176 60000
rect 50624 59600 50680 60000
rect 51128 59600 51184 60000
rect 51632 59600 51688 60000
rect 52136 59600 52192 60000
rect 52640 59600 52696 60000
rect 53144 59600 53200 60000
rect 53648 59600 53704 60000
rect 54152 59600 54208 60000
rect 54656 59600 54712 60000
rect 55160 59600 55216 60000
rect 55664 59600 55720 60000
rect 56168 59600 56224 60000
rect 56672 59600 56728 60000
rect 57176 59600 57232 60000
rect 57680 59600 57736 60000
rect 58184 59600 58240 60000
rect 58688 59600 58744 60000
rect 4984 0 5040 400
rect 5152 0 5208 400
rect 5320 0 5376 400
rect 5488 0 5544 400
rect 5656 0 5712 400
rect 5824 0 5880 400
rect 5992 0 6048 400
rect 6160 0 6216 400
rect 6328 0 6384 400
rect 6496 0 6552 400
rect 6664 0 6720 400
rect 6832 0 6888 400
rect 7000 0 7056 400
rect 7168 0 7224 400
rect 7336 0 7392 400
rect 7504 0 7560 400
rect 7672 0 7728 400
rect 7840 0 7896 400
rect 8008 0 8064 400
rect 8176 0 8232 400
rect 8344 0 8400 400
rect 8512 0 8568 400
rect 8680 0 8736 400
rect 8848 0 8904 400
rect 9016 0 9072 400
rect 9184 0 9240 400
rect 9352 0 9408 400
rect 9520 0 9576 400
rect 9688 0 9744 400
rect 9856 0 9912 400
rect 10024 0 10080 400
rect 10192 0 10248 400
rect 10360 0 10416 400
rect 10528 0 10584 400
rect 10696 0 10752 400
rect 10864 0 10920 400
rect 11032 0 11088 400
rect 11200 0 11256 400
rect 11368 0 11424 400
rect 11536 0 11592 400
rect 11704 0 11760 400
rect 11872 0 11928 400
rect 12040 0 12096 400
rect 12208 0 12264 400
rect 12376 0 12432 400
rect 12544 0 12600 400
rect 12712 0 12768 400
rect 12880 0 12936 400
rect 13048 0 13104 400
rect 13216 0 13272 400
rect 13384 0 13440 400
rect 13552 0 13608 400
rect 13720 0 13776 400
rect 13888 0 13944 400
rect 14056 0 14112 400
rect 14224 0 14280 400
rect 14392 0 14448 400
rect 14560 0 14616 400
rect 14728 0 14784 400
rect 14896 0 14952 400
rect 15064 0 15120 400
rect 15232 0 15288 400
rect 15400 0 15456 400
rect 15568 0 15624 400
rect 15736 0 15792 400
rect 15904 0 15960 400
rect 16072 0 16128 400
rect 16240 0 16296 400
rect 16408 0 16464 400
rect 16576 0 16632 400
rect 16744 0 16800 400
rect 16912 0 16968 400
rect 17080 0 17136 400
rect 17248 0 17304 400
rect 17416 0 17472 400
rect 17584 0 17640 400
rect 17752 0 17808 400
rect 17920 0 17976 400
rect 18088 0 18144 400
rect 18256 0 18312 400
rect 18424 0 18480 400
rect 18592 0 18648 400
rect 18760 0 18816 400
rect 18928 0 18984 400
rect 19096 0 19152 400
rect 19264 0 19320 400
rect 19432 0 19488 400
rect 19600 0 19656 400
rect 19768 0 19824 400
rect 19936 0 19992 400
rect 20104 0 20160 400
rect 20272 0 20328 400
rect 20440 0 20496 400
rect 20608 0 20664 400
rect 20776 0 20832 400
rect 20944 0 21000 400
rect 21112 0 21168 400
rect 21280 0 21336 400
rect 21448 0 21504 400
rect 21616 0 21672 400
rect 21784 0 21840 400
rect 21952 0 22008 400
rect 22120 0 22176 400
rect 22288 0 22344 400
rect 22456 0 22512 400
rect 22624 0 22680 400
rect 22792 0 22848 400
rect 22960 0 23016 400
rect 23128 0 23184 400
rect 23296 0 23352 400
rect 23464 0 23520 400
rect 23632 0 23688 400
rect 23800 0 23856 400
rect 23968 0 24024 400
rect 24136 0 24192 400
rect 24304 0 24360 400
rect 24472 0 24528 400
rect 24640 0 24696 400
rect 24808 0 24864 400
rect 24976 0 25032 400
rect 25144 0 25200 400
rect 25312 0 25368 400
rect 25480 0 25536 400
rect 25648 0 25704 400
rect 25816 0 25872 400
rect 25984 0 26040 400
rect 26152 0 26208 400
rect 26320 0 26376 400
rect 26488 0 26544 400
rect 26656 0 26712 400
rect 26824 0 26880 400
rect 26992 0 27048 400
rect 27160 0 27216 400
rect 27328 0 27384 400
rect 27496 0 27552 400
rect 27664 0 27720 400
rect 27832 0 27888 400
rect 28000 0 28056 400
rect 28168 0 28224 400
rect 28336 0 28392 400
rect 28504 0 28560 400
rect 28672 0 28728 400
rect 28840 0 28896 400
rect 29008 0 29064 400
rect 29176 0 29232 400
rect 29344 0 29400 400
rect 29512 0 29568 400
rect 29680 0 29736 400
rect 29848 0 29904 400
rect 30016 0 30072 400
rect 30184 0 30240 400
rect 30352 0 30408 400
rect 30520 0 30576 400
rect 30688 0 30744 400
rect 30856 0 30912 400
rect 31024 0 31080 400
rect 31192 0 31248 400
rect 31360 0 31416 400
rect 31528 0 31584 400
rect 31696 0 31752 400
rect 31864 0 31920 400
rect 32032 0 32088 400
rect 32200 0 32256 400
rect 32368 0 32424 400
rect 32536 0 32592 400
rect 32704 0 32760 400
rect 32872 0 32928 400
rect 33040 0 33096 400
rect 33208 0 33264 400
rect 33376 0 33432 400
rect 33544 0 33600 400
rect 33712 0 33768 400
rect 33880 0 33936 400
rect 34048 0 34104 400
rect 34216 0 34272 400
rect 34384 0 34440 400
rect 34552 0 34608 400
rect 34720 0 34776 400
rect 34888 0 34944 400
rect 35056 0 35112 400
rect 35224 0 35280 400
rect 35392 0 35448 400
rect 35560 0 35616 400
rect 35728 0 35784 400
rect 35896 0 35952 400
rect 36064 0 36120 400
rect 36232 0 36288 400
rect 36400 0 36456 400
rect 36568 0 36624 400
rect 36736 0 36792 400
rect 36904 0 36960 400
rect 37072 0 37128 400
rect 37240 0 37296 400
rect 37408 0 37464 400
rect 37576 0 37632 400
rect 37744 0 37800 400
rect 37912 0 37968 400
rect 38080 0 38136 400
rect 38248 0 38304 400
rect 38416 0 38472 400
rect 38584 0 38640 400
rect 38752 0 38808 400
rect 38920 0 38976 400
rect 39088 0 39144 400
rect 39256 0 39312 400
rect 39424 0 39480 400
rect 39592 0 39648 400
rect 39760 0 39816 400
rect 39928 0 39984 400
rect 40096 0 40152 400
rect 40264 0 40320 400
rect 40432 0 40488 400
rect 40600 0 40656 400
rect 40768 0 40824 400
rect 40936 0 40992 400
rect 41104 0 41160 400
rect 41272 0 41328 400
rect 41440 0 41496 400
rect 41608 0 41664 400
rect 41776 0 41832 400
rect 41944 0 42000 400
rect 42112 0 42168 400
rect 42280 0 42336 400
rect 42448 0 42504 400
rect 42616 0 42672 400
rect 42784 0 42840 400
rect 42952 0 43008 400
rect 43120 0 43176 400
rect 43288 0 43344 400
rect 43456 0 43512 400
rect 43624 0 43680 400
rect 43792 0 43848 400
rect 43960 0 44016 400
rect 44128 0 44184 400
rect 44296 0 44352 400
rect 44464 0 44520 400
rect 44632 0 44688 400
rect 44800 0 44856 400
rect 44968 0 45024 400
rect 45136 0 45192 400
rect 45304 0 45360 400
rect 45472 0 45528 400
rect 45640 0 45696 400
rect 45808 0 45864 400
rect 45976 0 46032 400
rect 46144 0 46200 400
rect 46312 0 46368 400
rect 46480 0 46536 400
rect 46648 0 46704 400
rect 46816 0 46872 400
rect 46984 0 47040 400
rect 47152 0 47208 400
rect 47320 0 47376 400
rect 47488 0 47544 400
rect 47656 0 47712 400
rect 47824 0 47880 400
rect 47992 0 48048 400
rect 48160 0 48216 400
rect 48328 0 48384 400
rect 48496 0 48552 400
rect 48664 0 48720 400
rect 48832 0 48888 400
rect 49000 0 49056 400
rect 49168 0 49224 400
rect 49336 0 49392 400
rect 49504 0 49560 400
rect 49672 0 49728 400
rect 49840 0 49896 400
rect 50008 0 50064 400
rect 50176 0 50232 400
rect 50344 0 50400 400
rect 50512 0 50568 400
rect 50680 0 50736 400
rect 50848 0 50904 400
rect 51016 0 51072 400
rect 51184 0 51240 400
rect 51352 0 51408 400
rect 51520 0 51576 400
rect 51688 0 51744 400
rect 51856 0 51912 400
rect 52024 0 52080 400
rect 52192 0 52248 400
rect 52360 0 52416 400
rect 52528 0 52584 400
rect 52696 0 52752 400
rect 52864 0 52920 400
rect 53032 0 53088 400
rect 53200 0 53256 400
rect 53368 0 53424 400
rect 53536 0 53592 400
rect 53704 0 53760 400
rect 53872 0 53928 400
rect 54040 0 54096 400
rect 54208 0 54264 400
rect 54376 0 54432 400
rect 54544 0 54600 400
rect 54712 0 54768 400
rect 54880 0 54936 400
<< obsm2 >>
rect 1134 59570 1202 59682
rect 1318 59570 1706 59682
rect 1822 59570 2210 59682
rect 2326 59570 2714 59682
rect 2830 59570 3218 59682
rect 3334 59570 3722 59682
rect 3838 59570 4226 59682
rect 4342 59570 4730 59682
rect 4846 59570 5234 59682
rect 5350 59570 5738 59682
rect 5854 59570 6242 59682
rect 6358 59570 6746 59682
rect 6862 59570 7250 59682
rect 7366 59570 7754 59682
rect 7870 59570 8258 59682
rect 8374 59570 8762 59682
rect 8878 59570 9266 59682
rect 9382 59570 9770 59682
rect 9886 59570 10274 59682
rect 10390 59570 10778 59682
rect 10894 59570 11282 59682
rect 11398 59570 11786 59682
rect 11902 59570 12290 59682
rect 12406 59570 12794 59682
rect 12910 59570 13298 59682
rect 13414 59570 13802 59682
rect 13918 59570 14306 59682
rect 14422 59570 14810 59682
rect 14926 59570 15314 59682
rect 15430 59570 15818 59682
rect 15934 59570 16322 59682
rect 16438 59570 16826 59682
rect 16942 59570 17330 59682
rect 17446 59570 17834 59682
rect 17950 59570 18338 59682
rect 18454 59570 18842 59682
rect 18958 59570 19346 59682
rect 19462 59570 19850 59682
rect 19966 59570 20354 59682
rect 20470 59570 20858 59682
rect 20974 59570 21362 59682
rect 21478 59570 21866 59682
rect 21982 59570 22370 59682
rect 22486 59570 22874 59682
rect 22990 59570 23378 59682
rect 23494 59570 23882 59682
rect 23998 59570 24386 59682
rect 24502 59570 24890 59682
rect 25006 59570 25394 59682
rect 25510 59570 25898 59682
rect 26014 59570 26402 59682
rect 26518 59570 26906 59682
rect 27022 59570 27410 59682
rect 27526 59570 27914 59682
rect 28030 59570 28418 59682
rect 28534 59570 28922 59682
rect 29038 59570 29426 59682
rect 29542 59570 29930 59682
rect 30046 59570 30434 59682
rect 30550 59570 30938 59682
rect 31054 59570 31442 59682
rect 31558 59570 31946 59682
rect 32062 59570 32450 59682
rect 32566 59570 32954 59682
rect 33070 59570 33458 59682
rect 33574 59570 33962 59682
rect 34078 59570 34466 59682
rect 34582 59570 34970 59682
rect 35086 59570 35474 59682
rect 35590 59570 35978 59682
rect 36094 59570 36482 59682
rect 36598 59570 36986 59682
rect 37102 59570 37490 59682
rect 37606 59570 37994 59682
rect 38110 59570 38498 59682
rect 38614 59570 39002 59682
rect 39118 59570 39506 59682
rect 39622 59570 40010 59682
rect 40126 59570 40514 59682
rect 40630 59570 41018 59682
rect 41134 59570 41522 59682
rect 41638 59570 42026 59682
rect 42142 59570 42530 59682
rect 42646 59570 43034 59682
rect 43150 59570 43538 59682
rect 43654 59570 44042 59682
rect 44158 59570 44546 59682
rect 44662 59570 45050 59682
rect 45166 59570 45554 59682
rect 45670 59570 46058 59682
rect 46174 59570 46562 59682
rect 46678 59570 47066 59682
rect 47182 59570 47570 59682
rect 47686 59570 48074 59682
rect 48190 59570 48578 59682
rect 48694 59570 49082 59682
rect 49198 59570 49586 59682
rect 49702 59570 50090 59682
rect 50206 59570 50594 59682
rect 50710 59570 51098 59682
rect 51214 59570 51602 59682
rect 51718 59570 52106 59682
rect 52222 59570 52610 59682
rect 52726 59570 53114 59682
rect 53230 59570 53618 59682
rect 53734 59570 54122 59682
rect 54238 59570 54626 59682
rect 54742 59570 55130 59682
rect 55246 59570 55634 59682
rect 55750 59570 56138 59682
rect 56254 59570 56642 59682
rect 56758 59570 57146 59682
rect 57262 59570 57650 59682
rect 57766 59570 58154 59682
rect 58270 59570 58658 59682
rect 58774 59570 58842 59682
rect 1134 430 58842 59570
rect 1134 400 4954 430
rect 5070 400 5122 430
rect 5238 400 5290 430
rect 5406 400 5458 430
rect 5574 400 5626 430
rect 5742 400 5794 430
rect 5910 400 5962 430
rect 6078 400 6130 430
rect 6246 400 6298 430
rect 6414 400 6466 430
rect 6582 400 6634 430
rect 6750 400 6802 430
rect 6918 400 6970 430
rect 7086 400 7138 430
rect 7254 400 7306 430
rect 7422 400 7474 430
rect 7590 400 7642 430
rect 7758 400 7810 430
rect 7926 400 7978 430
rect 8094 400 8146 430
rect 8262 400 8314 430
rect 8430 400 8482 430
rect 8598 400 8650 430
rect 8766 400 8818 430
rect 8934 400 8986 430
rect 9102 400 9154 430
rect 9270 400 9322 430
rect 9438 400 9490 430
rect 9606 400 9658 430
rect 9774 400 9826 430
rect 9942 400 9994 430
rect 10110 400 10162 430
rect 10278 400 10330 430
rect 10446 400 10498 430
rect 10614 400 10666 430
rect 10782 400 10834 430
rect 10950 400 11002 430
rect 11118 400 11170 430
rect 11286 400 11338 430
rect 11454 400 11506 430
rect 11622 400 11674 430
rect 11790 400 11842 430
rect 11958 400 12010 430
rect 12126 400 12178 430
rect 12294 400 12346 430
rect 12462 400 12514 430
rect 12630 400 12682 430
rect 12798 400 12850 430
rect 12966 400 13018 430
rect 13134 400 13186 430
rect 13302 400 13354 430
rect 13470 400 13522 430
rect 13638 400 13690 430
rect 13806 400 13858 430
rect 13974 400 14026 430
rect 14142 400 14194 430
rect 14310 400 14362 430
rect 14478 400 14530 430
rect 14646 400 14698 430
rect 14814 400 14866 430
rect 14982 400 15034 430
rect 15150 400 15202 430
rect 15318 400 15370 430
rect 15486 400 15538 430
rect 15654 400 15706 430
rect 15822 400 15874 430
rect 15990 400 16042 430
rect 16158 400 16210 430
rect 16326 400 16378 430
rect 16494 400 16546 430
rect 16662 400 16714 430
rect 16830 400 16882 430
rect 16998 400 17050 430
rect 17166 400 17218 430
rect 17334 400 17386 430
rect 17502 400 17554 430
rect 17670 400 17722 430
rect 17838 400 17890 430
rect 18006 400 18058 430
rect 18174 400 18226 430
rect 18342 400 18394 430
rect 18510 400 18562 430
rect 18678 400 18730 430
rect 18846 400 18898 430
rect 19014 400 19066 430
rect 19182 400 19234 430
rect 19350 400 19402 430
rect 19518 400 19570 430
rect 19686 400 19738 430
rect 19854 400 19906 430
rect 20022 400 20074 430
rect 20190 400 20242 430
rect 20358 400 20410 430
rect 20526 400 20578 430
rect 20694 400 20746 430
rect 20862 400 20914 430
rect 21030 400 21082 430
rect 21198 400 21250 430
rect 21366 400 21418 430
rect 21534 400 21586 430
rect 21702 400 21754 430
rect 21870 400 21922 430
rect 22038 400 22090 430
rect 22206 400 22258 430
rect 22374 400 22426 430
rect 22542 400 22594 430
rect 22710 400 22762 430
rect 22878 400 22930 430
rect 23046 400 23098 430
rect 23214 400 23266 430
rect 23382 400 23434 430
rect 23550 400 23602 430
rect 23718 400 23770 430
rect 23886 400 23938 430
rect 24054 400 24106 430
rect 24222 400 24274 430
rect 24390 400 24442 430
rect 24558 400 24610 430
rect 24726 400 24778 430
rect 24894 400 24946 430
rect 25062 400 25114 430
rect 25230 400 25282 430
rect 25398 400 25450 430
rect 25566 400 25618 430
rect 25734 400 25786 430
rect 25902 400 25954 430
rect 26070 400 26122 430
rect 26238 400 26290 430
rect 26406 400 26458 430
rect 26574 400 26626 430
rect 26742 400 26794 430
rect 26910 400 26962 430
rect 27078 400 27130 430
rect 27246 400 27298 430
rect 27414 400 27466 430
rect 27582 400 27634 430
rect 27750 400 27802 430
rect 27918 400 27970 430
rect 28086 400 28138 430
rect 28254 400 28306 430
rect 28422 400 28474 430
rect 28590 400 28642 430
rect 28758 400 28810 430
rect 28926 400 28978 430
rect 29094 400 29146 430
rect 29262 400 29314 430
rect 29430 400 29482 430
rect 29598 400 29650 430
rect 29766 400 29818 430
rect 29934 400 29986 430
rect 30102 400 30154 430
rect 30270 400 30322 430
rect 30438 400 30490 430
rect 30606 400 30658 430
rect 30774 400 30826 430
rect 30942 400 30994 430
rect 31110 400 31162 430
rect 31278 400 31330 430
rect 31446 400 31498 430
rect 31614 400 31666 430
rect 31782 400 31834 430
rect 31950 400 32002 430
rect 32118 400 32170 430
rect 32286 400 32338 430
rect 32454 400 32506 430
rect 32622 400 32674 430
rect 32790 400 32842 430
rect 32958 400 33010 430
rect 33126 400 33178 430
rect 33294 400 33346 430
rect 33462 400 33514 430
rect 33630 400 33682 430
rect 33798 400 33850 430
rect 33966 400 34018 430
rect 34134 400 34186 430
rect 34302 400 34354 430
rect 34470 400 34522 430
rect 34638 400 34690 430
rect 34806 400 34858 430
rect 34974 400 35026 430
rect 35142 400 35194 430
rect 35310 400 35362 430
rect 35478 400 35530 430
rect 35646 400 35698 430
rect 35814 400 35866 430
rect 35982 400 36034 430
rect 36150 400 36202 430
rect 36318 400 36370 430
rect 36486 400 36538 430
rect 36654 400 36706 430
rect 36822 400 36874 430
rect 36990 400 37042 430
rect 37158 400 37210 430
rect 37326 400 37378 430
rect 37494 400 37546 430
rect 37662 400 37714 430
rect 37830 400 37882 430
rect 37998 400 38050 430
rect 38166 400 38218 430
rect 38334 400 38386 430
rect 38502 400 38554 430
rect 38670 400 38722 430
rect 38838 400 38890 430
rect 39006 400 39058 430
rect 39174 400 39226 430
rect 39342 400 39394 430
rect 39510 400 39562 430
rect 39678 400 39730 430
rect 39846 400 39898 430
rect 40014 400 40066 430
rect 40182 400 40234 430
rect 40350 400 40402 430
rect 40518 400 40570 430
rect 40686 400 40738 430
rect 40854 400 40906 430
rect 41022 400 41074 430
rect 41190 400 41242 430
rect 41358 400 41410 430
rect 41526 400 41578 430
rect 41694 400 41746 430
rect 41862 400 41914 430
rect 42030 400 42082 430
rect 42198 400 42250 430
rect 42366 400 42418 430
rect 42534 400 42586 430
rect 42702 400 42754 430
rect 42870 400 42922 430
rect 43038 400 43090 430
rect 43206 400 43258 430
rect 43374 400 43426 430
rect 43542 400 43594 430
rect 43710 400 43762 430
rect 43878 400 43930 430
rect 44046 400 44098 430
rect 44214 400 44266 430
rect 44382 400 44434 430
rect 44550 400 44602 430
rect 44718 400 44770 430
rect 44886 400 44938 430
rect 45054 400 45106 430
rect 45222 400 45274 430
rect 45390 400 45442 430
rect 45558 400 45610 430
rect 45726 400 45778 430
rect 45894 400 45946 430
rect 46062 400 46114 430
rect 46230 400 46282 430
rect 46398 400 46450 430
rect 46566 400 46618 430
rect 46734 400 46786 430
rect 46902 400 46954 430
rect 47070 400 47122 430
rect 47238 400 47290 430
rect 47406 400 47458 430
rect 47574 400 47626 430
rect 47742 400 47794 430
rect 47910 400 47962 430
rect 48078 400 48130 430
rect 48246 400 48298 430
rect 48414 400 48466 430
rect 48582 400 48634 430
rect 48750 400 48802 430
rect 48918 400 48970 430
rect 49086 400 49138 430
rect 49254 400 49306 430
rect 49422 400 49474 430
rect 49590 400 49642 430
rect 49758 400 49810 430
rect 49926 400 49978 430
rect 50094 400 50146 430
rect 50262 400 50314 430
rect 50430 400 50482 430
rect 50598 400 50650 430
rect 50766 400 50818 430
rect 50934 400 50986 430
rect 51102 400 51154 430
rect 51270 400 51322 430
rect 51438 400 51490 430
rect 51606 400 51658 430
rect 51774 400 51826 430
rect 51942 400 51994 430
rect 52110 400 52162 430
rect 52278 400 52330 430
rect 52446 400 52498 430
rect 52614 400 52666 430
rect 52782 400 52834 430
rect 52950 400 53002 430
rect 53118 400 53170 430
rect 53286 400 53338 430
rect 53454 400 53506 430
rect 53622 400 53674 430
rect 53790 400 53842 430
rect 53958 400 54010 430
rect 54126 400 54178 430
rect 54294 400 54346 430
rect 54462 400 54514 430
rect 54630 400 54682 430
rect 54798 400 54850 430
rect 54966 400 58842 430
<< obsm3 >>
rect 2081 854 57783 58842
<< metal4 >>
rect 2224 1538 2384 58438
rect 9904 1538 10064 58438
rect 17584 1538 17744 58438
rect 25264 1538 25424 58438
rect 32944 1538 33104 58438
rect 40624 1538 40784 58438
rect 48304 1538 48464 58438
rect 55984 1538 56144 58438
<< obsm4 >>
rect 22638 55113 25234 58231
rect 25454 55113 32914 58231
rect 33134 55113 39466 58231
<< labels >>
rlabel metal2 s 1232 59600 1288 60000 6 io_active
port 1 nsew signal input
rlabel metal2 s 1736 59600 1792 60000 6 io_in[0]
port 2 nsew signal input
rlabel metal2 s 16856 59600 16912 60000 6 io_in[10]
port 3 nsew signal input
rlabel metal2 s 18368 59600 18424 60000 6 io_in[11]
port 4 nsew signal input
rlabel metal2 s 19880 59600 19936 60000 6 io_in[12]
port 5 nsew signal input
rlabel metal2 s 21392 59600 21448 60000 6 io_in[13]
port 6 nsew signal input
rlabel metal2 s 22904 59600 22960 60000 6 io_in[14]
port 7 nsew signal input
rlabel metal2 s 24416 59600 24472 60000 6 io_in[15]
port 8 nsew signal input
rlabel metal2 s 25928 59600 25984 60000 6 io_in[16]
port 9 nsew signal input
rlabel metal2 s 27440 59600 27496 60000 6 io_in[17]
port 10 nsew signal input
rlabel metal2 s 28952 59600 29008 60000 6 io_in[18]
port 11 nsew signal input
rlabel metal2 s 30464 59600 30520 60000 6 io_in[19]
port 12 nsew signal input
rlabel metal2 s 3248 59600 3304 60000 6 io_in[1]
port 13 nsew signal input
rlabel metal2 s 31976 59600 32032 60000 6 io_in[20]
port 14 nsew signal input
rlabel metal2 s 33488 59600 33544 60000 6 io_in[21]
port 15 nsew signal input
rlabel metal2 s 35000 59600 35056 60000 6 io_in[22]
port 16 nsew signal input
rlabel metal2 s 36512 59600 36568 60000 6 io_in[23]
port 17 nsew signal input
rlabel metal2 s 38024 59600 38080 60000 6 io_in[24]
port 18 nsew signal input
rlabel metal2 s 39536 59600 39592 60000 6 io_in[25]
port 19 nsew signal input
rlabel metal2 s 41048 59600 41104 60000 6 io_in[26]
port 20 nsew signal input
rlabel metal2 s 42560 59600 42616 60000 6 io_in[27]
port 21 nsew signal input
rlabel metal2 s 44072 59600 44128 60000 6 io_in[28]
port 22 nsew signal input
rlabel metal2 s 45584 59600 45640 60000 6 io_in[29]
port 23 nsew signal input
rlabel metal2 s 4760 59600 4816 60000 6 io_in[2]
port 24 nsew signal input
rlabel metal2 s 47096 59600 47152 60000 6 io_in[30]
port 25 nsew signal input
rlabel metal2 s 48608 59600 48664 60000 6 io_in[31]
port 26 nsew signal input
rlabel metal2 s 50120 59600 50176 60000 6 io_in[32]
port 27 nsew signal input
rlabel metal2 s 51632 59600 51688 60000 6 io_in[33]
port 28 nsew signal input
rlabel metal2 s 53144 59600 53200 60000 6 io_in[34]
port 29 nsew signal input
rlabel metal2 s 54656 59600 54712 60000 6 io_in[35]
port 30 nsew signal input
rlabel metal2 s 56168 59600 56224 60000 6 io_in[36]
port 31 nsew signal input
rlabel metal2 s 57680 59600 57736 60000 6 io_in[37]
port 32 nsew signal input
rlabel metal2 s 6272 59600 6328 60000 6 io_in[3]
port 33 nsew signal input
rlabel metal2 s 7784 59600 7840 60000 6 io_in[4]
port 34 nsew signal input
rlabel metal2 s 9296 59600 9352 60000 6 io_in[5]
port 35 nsew signal input
rlabel metal2 s 10808 59600 10864 60000 6 io_in[6]
port 36 nsew signal input
rlabel metal2 s 12320 59600 12376 60000 6 io_in[7]
port 37 nsew signal input
rlabel metal2 s 13832 59600 13888 60000 6 io_in[8]
port 38 nsew signal input
rlabel metal2 s 15344 59600 15400 60000 6 io_in[9]
port 39 nsew signal input
rlabel metal2 s 2240 59600 2296 60000 6 io_oeb[0]
port 40 nsew signal output
rlabel metal2 s 17360 59600 17416 60000 6 io_oeb[10]
port 41 nsew signal output
rlabel metal2 s 18872 59600 18928 60000 6 io_oeb[11]
port 42 nsew signal output
rlabel metal2 s 20384 59600 20440 60000 6 io_oeb[12]
port 43 nsew signal output
rlabel metal2 s 21896 59600 21952 60000 6 io_oeb[13]
port 44 nsew signal output
rlabel metal2 s 23408 59600 23464 60000 6 io_oeb[14]
port 45 nsew signal output
rlabel metal2 s 24920 59600 24976 60000 6 io_oeb[15]
port 46 nsew signal output
rlabel metal2 s 26432 59600 26488 60000 6 io_oeb[16]
port 47 nsew signal output
rlabel metal2 s 27944 59600 28000 60000 6 io_oeb[17]
port 48 nsew signal output
rlabel metal2 s 29456 59600 29512 60000 6 io_oeb[18]
port 49 nsew signal output
rlabel metal2 s 30968 59600 31024 60000 6 io_oeb[19]
port 50 nsew signal output
rlabel metal2 s 3752 59600 3808 60000 6 io_oeb[1]
port 51 nsew signal output
rlabel metal2 s 32480 59600 32536 60000 6 io_oeb[20]
port 52 nsew signal output
rlabel metal2 s 33992 59600 34048 60000 6 io_oeb[21]
port 53 nsew signal output
rlabel metal2 s 35504 59600 35560 60000 6 io_oeb[22]
port 54 nsew signal output
rlabel metal2 s 37016 59600 37072 60000 6 io_oeb[23]
port 55 nsew signal output
rlabel metal2 s 38528 59600 38584 60000 6 io_oeb[24]
port 56 nsew signal output
rlabel metal2 s 40040 59600 40096 60000 6 io_oeb[25]
port 57 nsew signal output
rlabel metal2 s 41552 59600 41608 60000 6 io_oeb[26]
port 58 nsew signal output
rlabel metal2 s 43064 59600 43120 60000 6 io_oeb[27]
port 59 nsew signal output
rlabel metal2 s 44576 59600 44632 60000 6 io_oeb[28]
port 60 nsew signal output
rlabel metal2 s 46088 59600 46144 60000 6 io_oeb[29]
port 61 nsew signal output
rlabel metal2 s 5264 59600 5320 60000 6 io_oeb[2]
port 62 nsew signal output
rlabel metal2 s 47600 59600 47656 60000 6 io_oeb[30]
port 63 nsew signal output
rlabel metal2 s 49112 59600 49168 60000 6 io_oeb[31]
port 64 nsew signal output
rlabel metal2 s 50624 59600 50680 60000 6 io_oeb[32]
port 65 nsew signal output
rlabel metal2 s 52136 59600 52192 60000 6 io_oeb[33]
port 66 nsew signal output
rlabel metal2 s 53648 59600 53704 60000 6 io_oeb[34]
port 67 nsew signal output
rlabel metal2 s 55160 59600 55216 60000 6 io_oeb[35]
port 68 nsew signal output
rlabel metal2 s 56672 59600 56728 60000 6 io_oeb[36]
port 69 nsew signal output
rlabel metal2 s 58184 59600 58240 60000 6 io_oeb[37]
port 70 nsew signal output
rlabel metal2 s 6776 59600 6832 60000 6 io_oeb[3]
port 71 nsew signal output
rlabel metal2 s 8288 59600 8344 60000 6 io_oeb[4]
port 72 nsew signal output
rlabel metal2 s 9800 59600 9856 60000 6 io_oeb[5]
port 73 nsew signal output
rlabel metal2 s 11312 59600 11368 60000 6 io_oeb[6]
port 74 nsew signal output
rlabel metal2 s 12824 59600 12880 60000 6 io_oeb[7]
port 75 nsew signal output
rlabel metal2 s 14336 59600 14392 60000 6 io_oeb[8]
port 76 nsew signal output
rlabel metal2 s 15848 59600 15904 60000 6 io_oeb[9]
port 77 nsew signal output
rlabel metal2 s 2744 59600 2800 60000 6 io_out[0]
port 78 nsew signal output
rlabel metal2 s 17864 59600 17920 60000 6 io_out[10]
port 79 nsew signal output
rlabel metal2 s 19376 59600 19432 60000 6 io_out[11]
port 80 nsew signal output
rlabel metal2 s 20888 59600 20944 60000 6 io_out[12]
port 81 nsew signal output
rlabel metal2 s 22400 59600 22456 60000 6 io_out[13]
port 82 nsew signal output
rlabel metal2 s 23912 59600 23968 60000 6 io_out[14]
port 83 nsew signal output
rlabel metal2 s 25424 59600 25480 60000 6 io_out[15]
port 84 nsew signal output
rlabel metal2 s 26936 59600 26992 60000 6 io_out[16]
port 85 nsew signal output
rlabel metal2 s 28448 59600 28504 60000 6 io_out[17]
port 86 nsew signal output
rlabel metal2 s 29960 59600 30016 60000 6 io_out[18]
port 87 nsew signal output
rlabel metal2 s 31472 59600 31528 60000 6 io_out[19]
port 88 nsew signal output
rlabel metal2 s 4256 59600 4312 60000 6 io_out[1]
port 89 nsew signal output
rlabel metal2 s 32984 59600 33040 60000 6 io_out[20]
port 90 nsew signal output
rlabel metal2 s 34496 59600 34552 60000 6 io_out[21]
port 91 nsew signal output
rlabel metal2 s 36008 59600 36064 60000 6 io_out[22]
port 92 nsew signal output
rlabel metal2 s 37520 59600 37576 60000 6 io_out[23]
port 93 nsew signal output
rlabel metal2 s 39032 59600 39088 60000 6 io_out[24]
port 94 nsew signal output
rlabel metal2 s 40544 59600 40600 60000 6 io_out[25]
port 95 nsew signal output
rlabel metal2 s 42056 59600 42112 60000 6 io_out[26]
port 96 nsew signal output
rlabel metal2 s 43568 59600 43624 60000 6 io_out[27]
port 97 nsew signal output
rlabel metal2 s 45080 59600 45136 60000 6 io_out[28]
port 98 nsew signal output
rlabel metal2 s 46592 59600 46648 60000 6 io_out[29]
port 99 nsew signal output
rlabel metal2 s 5768 59600 5824 60000 6 io_out[2]
port 100 nsew signal output
rlabel metal2 s 48104 59600 48160 60000 6 io_out[30]
port 101 nsew signal output
rlabel metal2 s 49616 59600 49672 60000 6 io_out[31]
port 102 nsew signal output
rlabel metal2 s 51128 59600 51184 60000 6 io_out[32]
port 103 nsew signal output
rlabel metal2 s 52640 59600 52696 60000 6 io_out[33]
port 104 nsew signal output
rlabel metal2 s 54152 59600 54208 60000 6 io_out[34]
port 105 nsew signal output
rlabel metal2 s 55664 59600 55720 60000 6 io_out[35]
port 106 nsew signal output
rlabel metal2 s 57176 59600 57232 60000 6 io_out[36]
port 107 nsew signal output
rlabel metal2 s 58688 59600 58744 60000 6 io_out[37]
port 108 nsew signal output
rlabel metal2 s 7280 59600 7336 60000 6 io_out[3]
port 109 nsew signal output
rlabel metal2 s 8792 59600 8848 60000 6 io_out[4]
port 110 nsew signal output
rlabel metal2 s 10304 59600 10360 60000 6 io_out[5]
port 111 nsew signal output
rlabel metal2 s 11816 59600 11872 60000 6 io_out[6]
port 112 nsew signal output
rlabel metal2 s 13328 59600 13384 60000 6 io_out[7]
port 113 nsew signal output
rlabel metal2 s 14840 59600 14896 60000 6 io_out[8]
port 114 nsew signal output
rlabel metal2 s 16352 59600 16408 60000 6 io_out[9]
port 115 nsew signal output
rlabel metal2 s 22792 0 22848 400 6 la_data_in[0]
port 116 nsew signal input
rlabel metal2 s 27832 0 27888 400 6 la_data_in[10]
port 117 nsew signal input
rlabel metal2 s 28336 0 28392 400 6 la_data_in[11]
port 118 nsew signal input
rlabel metal2 s 28840 0 28896 400 6 la_data_in[12]
port 119 nsew signal input
rlabel metal2 s 29344 0 29400 400 6 la_data_in[13]
port 120 nsew signal input
rlabel metal2 s 29848 0 29904 400 6 la_data_in[14]
port 121 nsew signal input
rlabel metal2 s 30352 0 30408 400 6 la_data_in[15]
port 122 nsew signal input
rlabel metal2 s 30856 0 30912 400 6 la_data_in[16]
port 123 nsew signal input
rlabel metal2 s 31360 0 31416 400 6 la_data_in[17]
port 124 nsew signal input
rlabel metal2 s 31864 0 31920 400 6 la_data_in[18]
port 125 nsew signal input
rlabel metal2 s 32368 0 32424 400 6 la_data_in[19]
port 126 nsew signal input
rlabel metal2 s 23296 0 23352 400 6 la_data_in[1]
port 127 nsew signal input
rlabel metal2 s 32872 0 32928 400 6 la_data_in[20]
port 128 nsew signal input
rlabel metal2 s 33376 0 33432 400 6 la_data_in[21]
port 129 nsew signal input
rlabel metal2 s 33880 0 33936 400 6 la_data_in[22]
port 130 nsew signal input
rlabel metal2 s 34384 0 34440 400 6 la_data_in[23]
port 131 nsew signal input
rlabel metal2 s 34888 0 34944 400 6 la_data_in[24]
port 132 nsew signal input
rlabel metal2 s 35392 0 35448 400 6 la_data_in[25]
port 133 nsew signal input
rlabel metal2 s 35896 0 35952 400 6 la_data_in[26]
port 134 nsew signal input
rlabel metal2 s 36400 0 36456 400 6 la_data_in[27]
port 135 nsew signal input
rlabel metal2 s 36904 0 36960 400 6 la_data_in[28]
port 136 nsew signal input
rlabel metal2 s 37408 0 37464 400 6 la_data_in[29]
port 137 nsew signal input
rlabel metal2 s 23800 0 23856 400 6 la_data_in[2]
port 138 nsew signal input
rlabel metal2 s 37912 0 37968 400 6 la_data_in[30]
port 139 nsew signal input
rlabel metal2 s 38416 0 38472 400 6 la_data_in[31]
port 140 nsew signal input
rlabel metal2 s 38920 0 38976 400 6 la_data_in[32]
port 141 nsew signal input
rlabel metal2 s 39424 0 39480 400 6 la_data_in[33]
port 142 nsew signal input
rlabel metal2 s 39928 0 39984 400 6 la_data_in[34]
port 143 nsew signal input
rlabel metal2 s 40432 0 40488 400 6 la_data_in[35]
port 144 nsew signal input
rlabel metal2 s 40936 0 40992 400 6 la_data_in[36]
port 145 nsew signal input
rlabel metal2 s 41440 0 41496 400 6 la_data_in[37]
port 146 nsew signal input
rlabel metal2 s 41944 0 42000 400 6 la_data_in[38]
port 147 nsew signal input
rlabel metal2 s 42448 0 42504 400 6 la_data_in[39]
port 148 nsew signal input
rlabel metal2 s 24304 0 24360 400 6 la_data_in[3]
port 149 nsew signal input
rlabel metal2 s 42952 0 43008 400 6 la_data_in[40]
port 150 nsew signal input
rlabel metal2 s 43456 0 43512 400 6 la_data_in[41]
port 151 nsew signal input
rlabel metal2 s 43960 0 44016 400 6 la_data_in[42]
port 152 nsew signal input
rlabel metal2 s 44464 0 44520 400 6 la_data_in[43]
port 153 nsew signal input
rlabel metal2 s 44968 0 45024 400 6 la_data_in[44]
port 154 nsew signal input
rlabel metal2 s 45472 0 45528 400 6 la_data_in[45]
port 155 nsew signal input
rlabel metal2 s 45976 0 46032 400 6 la_data_in[46]
port 156 nsew signal input
rlabel metal2 s 46480 0 46536 400 6 la_data_in[47]
port 157 nsew signal input
rlabel metal2 s 46984 0 47040 400 6 la_data_in[48]
port 158 nsew signal input
rlabel metal2 s 47488 0 47544 400 6 la_data_in[49]
port 159 nsew signal input
rlabel metal2 s 24808 0 24864 400 6 la_data_in[4]
port 160 nsew signal input
rlabel metal2 s 47992 0 48048 400 6 la_data_in[50]
port 161 nsew signal input
rlabel metal2 s 48496 0 48552 400 6 la_data_in[51]
port 162 nsew signal input
rlabel metal2 s 49000 0 49056 400 6 la_data_in[52]
port 163 nsew signal input
rlabel metal2 s 49504 0 49560 400 6 la_data_in[53]
port 164 nsew signal input
rlabel metal2 s 50008 0 50064 400 6 la_data_in[54]
port 165 nsew signal input
rlabel metal2 s 50512 0 50568 400 6 la_data_in[55]
port 166 nsew signal input
rlabel metal2 s 51016 0 51072 400 6 la_data_in[56]
port 167 nsew signal input
rlabel metal2 s 51520 0 51576 400 6 la_data_in[57]
port 168 nsew signal input
rlabel metal2 s 52024 0 52080 400 6 la_data_in[58]
port 169 nsew signal input
rlabel metal2 s 52528 0 52584 400 6 la_data_in[59]
port 170 nsew signal input
rlabel metal2 s 25312 0 25368 400 6 la_data_in[5]
port 171 nsew signal input
rlabel metal2 s 53032 0 53088 400 6 la_data_in[60]
port 172 nsew signal input
rlabel metal2 s 53536 0 53592 400 6 la_data_in[61]
port 173 nsew signal input
rlabel metal2 s 54040 0 54096 400 6 la_data_in[62]
port 174 nsew signal input
rlabel metal2 s 54544 0 54600 400 6 la_data_in[63]
port 175 nsew signal input
rlabel metal2 s 25816 0 25872 400 6 la_data_in[6]
port 176 nsew signal input
rlabel metal2 s 26320 0 26376 400 6 la_data_in[7]
port 177 nsew signal input
rlabel metal2 s 26824 0 26880 400 6 la_data_in[8]
port 178 nsew signal input
rlabel metal2 s 27328 0 27384 400 6 la_data_in[9]
port 179 nsew signal input
rlabel metal2 s 22960 0 23016 400 6 la_data_out[0]
port 180 nsew signal output
rlabel metal2 s 28000 0 28056 400 6 la_data_out[10]
port 181 nsew signal output
rlabel metal2 s 28504 0 28560 400 6 la_data_out[11]
port 182 nsew signal output
rlabel metal2 s 29008 0 29064 400 6 la_data_out[12]
port 183 nsew signal output
rlabel metal2 s 29512 0 29568 400 6 la_data_out[13]
port 184 nsew signal output
rlabel metal2 s 30016 0 30072 400 6 la_data_out[14]
port 185 nsew signal output
rlabel metal2 s 30520 0 30576 400 6 la_data_out[15]
port 186 nsew signal output
rlabel metal2 s 31024 0 31080 400 6 la_data_out[16]
port 187 nsew signal output
rlabel metal2 s 31528 0 31584 400 6 la_data_out[17]
port 188 nsew signal output
rlabel metal2 s 32032 0 32088 400 6 la_data_out[18]
port 189 nsew signal output
rlabel metal2 s 32536 0 32592 400 6 la_data_out[19]
port 190 nsew signal output
rlabel metal2 s 23464 0 23520 400 6 la_data_out[1]
port 191 nsew signal output
rlabel metal2 s 33040 0 33096 400 6 la_data_out[20]
port 192 nsew signal output
rlabel metal2 s 33544 0 33600 400 6 la_data_out[21]
port 193 nsew signal output
rlabel metal2 s 34048 0 34104 400 6 la_data_out[22]
port 194 nsew signal output
rlabel metal2 s 34552 0 34608 400 6 la_data_out[23]
port 195 nsew signal output
rlabel metal2 s 35056 0 35112 400 6 la_data_out[24]
port 196 nsew signal output
rlabel metal2 s 35560 0 35616 400 6 la_data_out[25]
port 197 nsew signal output
rlabel metal2 s 36064 0 36120 400 6 la_data_out[26]
port 198 nsew signal output
rlabel metal2 s 36568 0 36624 400 6 la_data_out[27]
port 199 nsew signal output
rlabel metal2 s 37072 0 37128 400 6 la_data_out[28]
port 200 nsew signal output
rlabel metal2 s 37576 0 37632 400 6 la_data_out[29]
port 201 nsew signal output
rlabel metal2 s 23968 0 24024 400 6 la_data_out[2]
port 202 nsew signal output
rlabel metal2 s 38080 0 38136 400 6 la_data_out[30]
port 203 nsew signal output
rlabel metal2 s 38584 0 38640 400 6 la_data_out[31]
port 204 nsew signal output
rlabel metal2 s 39088 0 39144 400 6 la_data_out[32]
port 205 nsew signal output
rlabel metal2 s 39592 0 39648 400 6 la_data_out[33]
port 206 nsew signal output
rlabel metal2 s 40096 0 40152 400 6 la_data_out[34]
port 207 nsew signal output
rlabel metal2 s 40600 0 40656 400 6 la_data_out[35]
port 208 nsew signal output
rlabel metal2 s 41104 0 41160 400 6 la_data_out[36]
port 209 nsew signal output
rlabel metal2 s 41608 0 41664 400 6 la_data_out[37]
port 210 nsew signal output
rlabel metal2 s 42112 0 42168 400 6 la_data_out[38]
port 211 nsew signal output
rlabel metal2 s 42616 0 42672 400 6 la_data_out[39]
port 212 nsew signal output
rlabel metal2 s 24472 0 24528 400 6 la_data_out[3]
port 213 nsew signal output
rlabel metal2 s 43120 0 43176 400 6 la_data_out[40]
port 214 nsew signal output
rlabel metal2 s 43624 0 43680 400 6 la_data_out[41]
port 215 nsew signal output
rlabel metal2 s 44128 0 44184 400 6 la_data_out[42]
port 216 nsew signal output
rlabel metal2 s 44632 0 44688 400 6 la_data_out[43]
port 217 nsew signal output
rlabel metal2 s 45136 0 45192 400 6 la_data_out[44]
port 218 nsew signal output
rlabel metal2 s 45640 0 45696 400 6 la_data_out[45]
port 219 nsew signal output
rlabel metal2 s 46144 0 46200 400 6 la_data_out[46]
port 220 nsew signal output
rlabel metal2 s 46648 0 46704 400 6 la_data_out[47]
port 221 nsew signal output
rlabel metal2 s 47152 0 47208 400 6 la_data_out[48]
port 222 nsew signal output
rlabel metal2 s 47656 0 47712 400 6 la_data_out[49]
port 223 nsew signal output
rlabel metal2 s 24976 0 25032 400 6 la_data_out[4]
port 224 nsew signal output
rlabel metal2 s 48160 0 48216 400 6 la_data_out[50]
port 225 nsew signal output
rlabel metal2 s 48664 0 48720 400 6 la_data_out[51]
port 226 nsew signal output
rlabel metal2 s 49168 0 49224 400 6 la_data_out[52]
port 227 nsew signal output
rlabel metal2 s 49672 0 49728 400 6 la_data_out[53]
port 228 nsew signal output
rlabel metal2 s 50176 0 50232 400 6 la_data_out[54]
port 229 nsew signal output
rlabel metal2 s 50680 0 50736 400 6 la_data_out[55]
port 230 nsew signal output
rlabel metal2 s 51184 0 51240 400 6 la_data_out[56]
port 231 nsew signal output
rlabel metal2 s 51688 0 51744 400 6 la_data_out[57]
port 232 nsew signal output
rlabel metal2 s 52192 0 52248 400 6 la_data_out[58]
port 233 nsew signal output
rlabel metal2 s 52696 0 52752 400 6 la_data_out[59]
port 234 nsew signal output
rlabel metal2 s 25480 0 25536 400 6 la_data_out[5]
port 235 nsew signal output
rlabel metal2 s 53200 0 53256 400 6 la_data_out[60]
port 236 nsew signal output
rlabel metal2 s 53704 0 53760 400 6 la_data_out[61]
port 237 nsew signal output
rlabel metal2 s 54208 0 54264 400 6 la_data_out[62]
port 238 nsew signal output
rlabel metal2 s 54712 0 54768 400 6 la_data_out[63]
port 239 nsew signal output
rlabel metal2 s 25984 0 26040 400 6 la_data_out[6]
port 240 nsew signal output
rlabel metal2 s 26488 0 26544 400 6 la_data_out[7]
port 241 nsew signal output
rlabel metal2 s 26992 0 27048 400 6 la_data_out[8]
port 242 nsew signal output
rlabel metal2 s 27496 0 27552 400 6 la_data_out[9]
port 243 nsew signal output
rlabel metal2 s 23128 0 23184 400 6 la_oenb[0]
port 244 nsew signal input
rlabel metal2 s 28168 0 28224 400 6 la_oenb[10]
port 245 nsew signal input
rlabel metal2 s 28672 0 28728 400 6 la_oenb[11]
port 246 nsew signal input
rlabel metal2 s 29176 0 29232 400 6 la_oenb[12]
port 247 nsew signal input
rlabel metal2 s 29680 0 29736 400 6 la_oenb[13]
port 248 nsew signal input
rlabel metal2 s 30184 0 30240 400 6 la_oenb[14]
port 249 nsew signal input
rlabel metal2 s 30688 0 30744 400 6 la_oenb[15]
port 250 nsew signal input
rlabel metal2 s 31192 0 31248 400 6 la_oenb[16]
port 251 nsew signal input
rlabel metal2 s 31696 0 31752 400 6 la_oenb[17]
port 252 nsew signal input
rlabel metal2 s 32200 0 32256 400 6 la_oenb[18]
port 253 nsew signal input
rlabel metal2 s 32704 0 32760 400 6 la_oenb[19]
port 254 nsew signal input
rlabel metal2 s 23632 0 23688 400 6 la_oenb[1]
port 255 nsew signal input
rlabel metal2 s 33208 0 33264 400 6 la_oenb[20]
port 256 nsew signal input
rlabel metal2 s 33712 0 33768 400 6 la_oenb[21]
port 257 nsew signal input
rlabel metal2 s 34216 0 34272 400 6 la_oenb[22]
port 258 nsew signal input
rlabel metal2 s 34720 0 34776 400 6 la_oenb[23]
port 259 nsew signal input
rlabel metal2 s 35224 0 35280 400 6 la_oenb[24]
port 260 nsew signal input
rlabel metal2 s 35728 0 35784 400 6 la_oenb[25]
port 261 nsew signal input
rlabel metal2 s 36232 0 36288 400 6 la_oenb[26]
port 262 nsew signal input
rlabel metal2 s 36736 0 36792 400 6 la_oenb[27]
port 263 nsew signal input
rlabel metal2 s 37240 0 37296 400 6 la_oenb[28]
port 264 nsew signal input
rlabel metal2 s 37744 0 37800 400 6 la_oenb[29]
port 265 nsew signal input
rlabel metal2 s 24136 0 24192 400 6 la_oenb[2]
port 266 nsew signal input
rlabel metal2 s 38248 0 38304 400 6 la_oenb[30]
port 267 nsew signal input
rlabel metal2 s 38752 0 38808 400 6 la_oenb[31]
port 268 nsew signal input
rlabel metal2 s 39256 0 39312 400 6 la_oenb[32]
port 269 nsew signal input
rlabel metal2 s 39760 0 39816 400 6 la_oenb[33]
port 270 nsew signal input
rlabel metal2 s 40264 0 40320 400 6 la_oenb[34]
port 271 nsew signal input
rlabel metal2 s 40768 0 40824 400 6 la_oenb[35]
port 272 nsew signal input
rlabel metal2 s 41272 0 41328 400 6 la_oenb[36]
port 273 nsew signal input
rlabel metal2 s 41776 0 41832 400 6 la_oenb[37]
port 274 nsew signal input
rlabel metal2 s 42280 0 42336 400 6 la_oenb[38]
port 275 nsew signal input
rlabel metal2 s 42784 0 42840 400 6 la_oenb[39]
port 276 nsew signal input
rlabel metal2 s 24640 0 24696 400 6 la_oenb[3]
port 277 nsew signal input
rlabel metal2 s 43288 0 43344 400 6 la_oenb[40]
port 278 nsew signal input
rlabel metal2 s 43792 0 43848 400 6 la_oenb[41]
port 279 nsew signal input
rlabel metal2 s 44296 0 44352 400 6 la_oenb[42]
port 280 nsew signal input
rlabel metal2 s 44800 0 44856 400 6 la_oenb[43]
port 281 nsew signal input
rlabel metal2 s 45304 0 45360 400 6 la_oenb[44]
port 282 nsew signal input
rlabel metal2 s 45808 0 45864 400 6 la_oenb[45]
port 283 nsew signal input
rlabel metal2 s 46312 0 46368 400 6 la_oenb[46]
port 284 nsew signal input
rlabel metal2 s 46816 0 46872 400 6 la_oenb[47]
port 285 nsew signal input
rlabel metal2 s 47320 0 47376 400 6 la_oenb[48]
port 286 nsew signal input
rlabel metal2 s 47824 0 47880 400 6 la_oenb[49]
port 287 nsew signal input
rlabel metal2 s 25144 0 25200 400 6 la_oenb[4]
port 288 nsew signal input
rlabel metal2 s 48328 0 48384 400 6 la_oenb[50]
port 289 nsew signal input
rlabel metal2 s 48832 0 48888 400 6 la_oenb[51]
port 290 nsew signal input
rlabel metal2 s 49336 0 49392 400 6 la_oenb[52]
port 291 nsew signal input
rlabel metal2 s 49840 0 49896 400 6 la_oenb[53]
port 292 nsew signal input
rlabel metal2 s 50344 0 50400 400 6 la_oenb[54]
port 293 nsew signal input
rlabel metal2 s 50848 0 50904 400 6 la_oenb[55]
port 294 nsew signal input
rlabel metal2 s 51352 0 51408 400 6 la_oenb[56]
port 295 nsew signal input
rlabel metal2 s 51856 0 51912 400 6 la_oenb[57]
port 296 nsew signal input
rlabel metal2 s 52360 0 52416 400 6 la_oenb[58]
port 297 nsew signal input
rlabel metal2 s 52864 0 52920 400 6 la_oenb[59]
port 298 nsew signal input
rlabel metal2 s 25648 0 25704 400 6 la_oenb[5]
port 299 nsew signal input
rlabel metal2 s 53368 0 53424 400 6 la_oenb[60]
port 300 nsew signal input
rlabel metal2 s 53872 0 53928 400 6 la_oenb[61]
port 301 nsew signal input
rlabel metal2 s 54376 0 54432 400 6 la_oenb[62]
port 302 nsew signal input
rlabel metal2 s 54880 0 54936 400 6 la_oenb[63]
port 303 nsew signal input
rlabel metal2 s 26152 0 26208 400 6 la_oenb[6]
port 304 nsew signal input
rlabel metal2 s 26656 0 26712 400 6 la_oenb[7]
port 305 nsew signal input
rlabel metal2 s 27160 0 27216 400 6 la_oenb[8]
port 306 nsew signal input
rlabel metal2 s 27664 0 27720 400 6 la_oenb[9]
port 307 nsew signal input
rlabel metal4 s 2224 1538 2384 58438 6 vdd
port 308 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 58438 6 vdd
port 308 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 58438 6 vdd
port 308 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 58438 6 vdd
port 308 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 58438 6 vss
port 309 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 58438 6 vss
port 309 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 58438 6 vss
port 309 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 58438 6 vss
port 309 nsew ground bidirectional
rlabel metal2 s 4984 0 5040 400 6 wb_clk_i
port 310 nsew signal input
rlabel metal2 s 5152 0 5208 400 6 wb_rst_i
port 311 nsew signal input
rlabel metal2 s 5320 0 5376 400 6 wbs_ack_o
port 312 nsew signal output
rlabel metal2 s 5992 0 6048 400 6 wbs_adr_i[0]
port 313 nsew signal input
rlabel metal2 s 11704 0 11760 400 6 wbs_adr_i[10]
port 314 nsew signal input
rlabel metal2 s 12208 0 12264 400 6 wbs_adr_i[11]
port 315 nsew signal input
rlabel metal2 s 12712 0 12768 400 6 wbs_adr_i[12]
port 316 nsew signal input
rlabel metal2 s 13216 0 13272 400 6 wbs_adr_i[13]
port 317 nsew signal input
rlabel metal2 s 13720 0 13776 400 6 wbs_adr_i[14]
port 318 nsew signal input
rlabel metal2 s 14224 0 14280 400 6 wbs_adr_i[15]
port 319 nsew signal input
rlabel metal2 s 14728 0 14784 400 6 wbs_adr_i[16]
port 320 nsew signal input
rlabel metal2 s 15232 0 15288 400 6 wbs_adr_i[17]
port 321 nsew signal input
rlabel metal2 s 15736 0 15792 400 6 wbs_adr_i[18]
port 322 nsew signal input
rlabel metal2 s 16240 0 16296 400 6 wbs_adr_i[19]
port 323 nsew signal input
rlabel metal2 s 6664 0 6720 400 6 wbs_adr_i[1]
port 324 nsew signal input
rlabel metal2 s 16744 0 16800 400 6 wbs_adr_i[20]
port 325 nsew signal input
rlabel metal2 s 17248 0 17304 400 6 wbs_adr_i[21]
port 326 nsew signal input
rlabel metal2 s 17752 0 17808 400 6 wbs_adr_i[22]
port 327 nsew signal input
rlabel metal2 s 18256 0 18312 400 6 wbs_adr_i[23]
port 328 nsew signal input
rlabel metal2 s 18760 0 18816 400 6 wbs_adr_i[24]
port 329 nsew signal input
rlabel metal2 s 19264 0 19320 400 6 wbs_adr_i[25]
port 330 nsew signal input
rlabel metal2 s 19768 0 19824 400 6 wbs_adr_i[26]
port 331 nsew signal input
rlabel metal2 s 20272 0 20328 400 6 wbs_adr_i[27]
port 332 nsew signal input
rlabel metal2 s 20776 0 20832 400 6 wbs_adr_i[28]
port 333 nsew signal input
rlabel metal2 s 21280 0 21336 400 6 wbs_adr_i[29]
port 334 nsew signal input
rlabel metal2 s 7336 0 7392 400 6 wbs_adr_i[2]
port 335 nsew signal input
rlabel metal2 s 21784 0 21840 400 6 wbs_adr_i[30]
port 336 nsew signal input
rlabel metal2 s 22288 0 22344 400 6 wbs_adr_i[31]
port 337 nsew signal input
rlabel metal2 s 8008 0 8064 400 6 wbs_adr_i[3]
port 338 nsew signal input
rlabel metal2 s 8680 0 8736 400 6 wbs_adr_i[4]
port 339 nsew signal input
rlabel metal2 s 9184 0 9240 400 6 wbs_adr_i[5]
port 340 nsew signal input
rlabel metal2 s 9688 0 9744 400 6 wbs_adr_i[6]
port 341 nsew signal input
rlabel metal2 s 10192 0 10248 400 6 wbs_adr_i[7]
port 342 nsew signal input
rlabel metal2 s 10696 0 10752 400 6 wbs_adr_i[8]
port 343 nsew signal input
rlabel metal2 s 11200 0 11256 400 6 wbs_adr_i[9]
port 344 nsew signal input
rlabel metal2 s 5488 0 5544 400 6 wbs_cyc_i
port 345 nsew signal input
rlabel metal2 s 6160 0 6216 400 6 wbs_dat_i[0]
port 346 nsew signal input
rlabel metal2 s 11872 0 11928 400 6 wbs_dat_i[10]
port 347 nsew signal input
rlabel metal2 s 12376 0 12432 400 6 wbs_dat_i[11]
port 348 nsew signal input
rlabel metal2 s 12880 0 12936 400 6 wbs_dat_i[12]
port 349 nsew signal input
rlabel metal2 s 13384 0 13440 400 6 wbs_dat_i[13]
port 350 nsew signal input
rlabel metal2 s 13888 0 13944 400 6 wbs_dat_i[14]
port 351 nsew signal input
rlabel metal2 s 14392 0 14448 400 6 wbs_dat_i[15]
port 352 nsew signal input
rlabel metal2 s 14896 0 14952 400 6 wbs_dat_i[16]
port 353 nsew signal input
rlabel metal2 s 15400 0 15456 400 6 wbs_dat_i[17]
port 354 nsew signal input
rlabel metal2 s 15904 0 15960 400 6 wbs_dat_i[18]
port 355 nsew signal input
rlabel metal2 s 16408 0 16464 400 6 wbs_dat_i[19]
port 356 nsew signal input
rlabel metal2 s 6832 0 6888 400 6 wbs_dat_i[1]
port 357 nsew signal input
rlabel metal2 s 16912 0 16968 400 6 wbs_dat_i[20]
port 358 nsew signal input
rlabel metal2 s 17416 0 17472 400 6 wbs_dat_i[21]
port 359 nsew signal input
rlabel metal2 s 17920 0 17976 400 6 wbs_dat_i[22]
port 360 nsew signal input
rlabel metal2 s 18424 0 18480 400 6 wbs_dat_i[23]
port 361 nsew signal input
rlabel metal2 s 18928 0 18984 400 6 wbs_dat_i[24]
port 362 nsew signal input
rlabel metal2 s 19432 0 19488 400 6 wbs_dat_i[25]
port 363 nsew signal input
rlabel metal2 s 19936 0 19992 400 6 wbs_dat_i[26]
port 364 nsew signal input
rlabel metal2 s 20440 0 20496 400 6 wbs_dat_i[27]
port 365 nsew signal input
rlabel metal2 s 20944 0 21000 400 6 wbs_dat_i[28]
port 366 nsew signal input
rlabel metal2 s 21448 0 21504 400 6 wbs_dat_i[29]
port 367 nsew signal input
rlabel metal2 s 7504 0 7560 400 6 wbs_dat_i[2]
port 368 nsew signal input
rlabel metal2 s 21952 0 22008 400 6 wbs_dat_i[30]
port 369 nsew signal input
rlabel metal2 s 22456 0 22512 400 6 wbs_dat_i[31]
port 370 nsew signal input
rlabel metal2 s 8176 0 8232 400 6 wbs_dat_i[3]
port 371 nsew signal input
rlabel metal2 s 8848 0 8904 400 6 wbs_dat_i[4]
port 372 nsew signal input
rlabel metal2 s 9352 0 9408 400 6 wbs_dat_i[5]
port 373 nsew signal input
rlabel metal2 s 9856 0 9912 400 6 wbs_dat_i[6]
port 374 nsew signal input
rlabel metal2 s 10360 0 10416 400 6 wbs_dat_i[7]
port 375 nsew signal input
rlabel metal2 s 10864 0 10920 400 6 wbs_dat_i[8]
port 376 nsew signal input
rlabel metal2 s 11368 0 11424 400 6 wbs_dat_i[9]
port 377 nsew signal input
rlabel metal2 s 6328 0 6384 400 6 wbs_dat_o[0]
port 378 nsew signal output
rlabel metal2 s 12040 0 12096 400 6 wbs_dat_o[10]
port 379 nsew signal output
rlabel metal2 s 12544 0 12600 400 6 wbs_dat_o[11]
port 380 nsew signal output
rlabel metal2 s 13048 0 13104 400 6 wbs_dat_o[12]
port 381 nsew signal output
rlabel metal2 s 13552 0 13608 400 6 wbs_dat_o[13]
port 382 nsew signal output
rlabel metal2 s 14056 0 14112 400 6 wbs_dat_o[14]
port 383 nsew signal output
rlabel metal2 s 14560 0 14616 400 6 wbs_dat_o[15]
port 384 nsew signal output
rlabel metal2 s 15064 0 15120 400 6 wbs_dat_o[16]
port 385 nsew signal output
rlabel metal2 s 15568 0 15624 400 6 wbs_dat_o[17]
port 386 nsew signal output
rlabel metal2 s 16072 0 16128 400 6 wbs_dat_o[18]
port 387 nsew signal output
rlabel metal2 s 16576 0 16632 400 6 wbs_dat_o[19]
port 388 nsew signal output
rlabel metal2 s 7000 0 7056 400 6 wbs_dat_o[1]
port 389 nsew signal output
rlabel metal2 s 17080 0 17136 400 6 wbs_dat_o[20]
port 390 nsew signal output
rlabel metal2 s 17584 0 17640 400 6 wbs_dat_o[21]
port 391 nsew signal output
rlabel metal2 s 18088 0 18144 400 6 wbs_dat_o[22]
port 392 nsew signal output
rlabel metal2 s 18592 0 18648 400 6 wbs_dat_o[23]
port 393 nsew signal output
rlabel metal2 s 19096 0 19152 400 6 wbs_dat_o[24]
port 394 nsew signal output
rlabel metal2 s 19600 0 19656 400 6 wbs_dat_o[25]
port 395 nsew signal output
rlabel metal2 s 20104 0 20160 400 6 wbs_dat_o[26]
port 396 nsew signal output
rlabel metal2 s 20608 0 20664 400 6 wbs_dat_o[27]
port 397 nsew signal output
rlabel metal2 s 21112 0 21168 400 6 wbs_dat_o[28]
port 398 nsew signal output
rlabel metal2 s 21616 0 21672 400 6 wbs_dat_o[29]
port 399 nsew signal output
rlabel metal2 s 7672 0 7728 400 6 wbs_dat_o[2]
port 400 nsew signal output
rlabel metal2 s 22120 0 22176 400 6 wbs_dat_o[30]
port 401 nsew signal output
rlabel metal2 s 22624 0 22680 400 6 wbs_dat_o[31]
port 402 nsew signal output
rlabel metal2 s 8344 0 8400 400 6 wbs_dat_o[3]
port 403 nsew signal output
rlabel metal2 s 9016 0 9072 400 6 wbs_dat_o[4]
port 404 nsew signal output
rlabel metal2 s 9520 0 9576 400 6 wbs_dat_o[5]
port 405 nsew signal output
rlabel metal2 s 10024 0 10080 400 6 wbs_dat_o[6]
port 406 nsew signal output
rlabel metal2 s 10528 0 10584 400 6 wbs_dat_o[7]
port 407 nsew signal output
rlabel metal2 s 11032 0 11088 400 6 wbs_dat_o[8]
port 408 nsew signal output
rlabel metal2 s 11536 0 11592 400 6 wbs_dat_o[9]
port 409 nsew signal output
rlabel metal2 s 6496 0 6552 400 6 wbs_sel_i[0]
port 410 nsew signal input
rlabel metal2 s 7168 0 7224 400 6 wbs_sel_i[1]
port 411 nsew signal input
rlabel metal2 s 7840 0 7896 400 6 wbs_sel_i[2]
port 412 nsew signal input
rlabel metal2 s 8512 0 8568 400 6 wbs_sel_i[3]
port 413 nsew signal input
rlabel metal2 s 5656 0 5712 400 6 wbs_stb_i
port 414 nsew signal input
rlabel metal2 s 5824 0 5880 400 6 wbs_we_i
port 415 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1835964
string GDS_FILE /opt/caravel_180/openlane/user_proj_example/runs/22_12_05_06_59/results/signoff/macro_golden.magic.gds
string GDS_START 162254
<< end >>

