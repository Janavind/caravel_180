VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2980.200 BY 2980.200 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 1209.320 2985.000 1210.440 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2271.640 2977.800 2272.760 2985.000 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1942.360 2977.800 1943.480 2985.000 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1613.080 2977.800 1614.200 2985.000 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1283.800 2977.800 1284.920 2985.000 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 954.520 2977.800 955.640 2985.000 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 625.240 2977.800 626.360 2985.000 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 295.960 2977.800 297.080 2985.000 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2943.640 2.400 2944.760 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2724.120 2.400 2725.240 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2504.600 2.400 2505.720 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 1433.320 2985.000 1434.440 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2285.080 2.400 2286.200 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2065.560 2.400 2066.680 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1846.040 2.400 1847.160 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1626.520 2.400 1627.640 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1407.000 2.400 1408.120 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1187.480 2.400 1188.600 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 967.960 2.400 969.080 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 748.440 2.400 749.560 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 528.920 2.400 530.040 ;
    END
  END analog_io[28]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 1657.320 2985.000 1658.440 ;
    END
  END analog_io[2]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 1881.320 2985.000 1882.440 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 2105.320 2985.000 2106.440 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 2329.320 2985.000 2330.440 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 2553.320 2985.000 2554.440 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 2777.320 2985.000 2778.440 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2930.200 2977.800 2931.320 2985.000 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2600.920 2977.800 2602.040 2985.000 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 33.320 2985.000 34.440 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 1937.320 2985.000 1938.440 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 2161.320 2985.000 2162.440 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 2385.320 2985.000 2386.440 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 2609.320 2985.000 2610.440 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 2833.320 2985.000 2834.440 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2847.880 2977.800 2849.000 2985.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2518.600 2977.800 2519.720 2985.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2189.320 2977.800 2190.440 2985.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1860.040 2977.800 1861.160 2985.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1530.760 2977.800 1531.880 2985.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 201.320 2985.000 202.440 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1201.480 2977.800 1202.600 2985.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 872.200 2977.800 873.320 2985.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 542.920 2977.800 544.040 2985.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 213.640 2977.800 214.760 2985.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2888.760 2.400 2889.880 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2669.240 2.400 2670.360 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2449.720 2.400 2450.840 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2230.200 2.400 2231.320 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2010.680 2.400 2011.800 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1791.160 2.400 1792.280 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 369.320 2985.000 370.440 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1571.640 2.400 1572.760 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1352.120 2.400 1353.240 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1132.600 2.400 1133.720 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 913.080 2.400 914.200 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 693.560 2.400 694.680 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 474.040 2.400 475.160 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 309.400 2.400 310.520 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 144.760 2.400 145.880 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 537.320 2985.000 538.440 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 705.320 2985.000 706.440 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 873.320 2985.000 874.440 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 1041.320 2985.000 1042.440 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 1265.320 2985.000 1266.440 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 1489.320 2985.000 1490.440 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 1713.320 2985.000 1714.440 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 145.320 2985.000 146.440 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 2049.320 2985.000 2050.440 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 2273.320 2985.000 2274.440 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 2497.320 2985.000 2498.440 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 2721.320 2985.000 2722.440 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 2945.320 2985.000 2946.440 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2683.240 2977.800 2684.360 2985.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2353.960 2977.800 2355.080 2985.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2024.680 2977.800 2025.800 2985.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1695.400 2977.800 1696.520 2985.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1366.120 2977.800 1367.240 2985.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 313.320 2985.000 314.440 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1036.840 2977.800 1037.960 2985.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 707.560 2977.800 708.680 2985.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 378.280 2977.800 379.400 2985.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 49.000 2977.800 50.120 2985.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2779.000 2.400 2780.120 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2559.480 2.400 2560.600 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2339.960 2.400 2341.080 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2120.440 2.400 2121.560 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1900.920 2.400 1902.040 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1681.400 2.400 1682.520 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 481.320 2985.000 482.440 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1461.880 2.400 1463.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1242.360 2.400 1243.480 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1022.840 2.400 1023.960 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 803.320 2.400 804.440 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 583.800 2.400 584.920 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 364.280 2.400 365.400 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 199.640 2.400 200.760 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 35.000 2.400 36.120 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 649.320 2985.000 650.440 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 817.320 2985.000 818.440 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 985.320 2985.000 986.440 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 1153.320 2985.000 1154.440 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 1377.320 2985.000 1378.440 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 1601.320 2985.000 1602.440 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 1825.320 2985.000 1826.440 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 89.320 2985.000 90.440 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 1993.320 2985.000 1994.440 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 2217.320 2985.000 2218.440 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 2441.320 2985.000 2442.440 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 2665.320 2985.000 2666.440 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 2889.320 2985.000 2890.440 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2765.560 2977.800 2766.680 2985.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2436.280 2977.800 2437.400 2985.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2107.000 2977.800 2108.120 2985.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1777.720 2977.800 1778.840 2985.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1448.440 2977.800 1449.560 2985.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 257.320 2985.000 258.440 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1119.160 2977.800 1120.280 2985.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 789.880 2977.800 791.000 2985.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 460.600 2977.800 461.720 2985.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 131.320 2977.800 132.440 2985.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2833.880 2.400 2835.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2614.360 2.400 2615.480 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2394.840 2.400 2395.960 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2175.320 2.400 2176.440 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1955.800 2.400 1956.920 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1736.280 2.400 1737.400 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 425.320 2985.000 426.440 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1516.760 2.400 1517.880 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1297.240 2.400 1298.360 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1077.720 2.400 1078.840 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 858.200 2.400 859.320 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 638.680 2.400 639.800 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 419.160 2.400 420.280 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 254.520 2.400 255.640 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 89.880 2.400 91.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 593.320 2985.000 594.440 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 761.320 2985.000 762.440 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 929.320 2985.000 930.440 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 1097.320 2985.000 1098.440 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 1321.320 2985.000 1322.440 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 1545.320 2985.000 1546.440 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2977.800 1769.320 2985.000 1770.440 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 702.520 -4.800 703.640 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2382.520 -4.800 2383.640 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2399.320 -4.800 2400.440 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2416.120 -4.800 2417.240 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2432.920 -4.800 2434.040 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2449.720 -4.800 2450.840 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2466.520 -4.800 2467.640 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2483.320 -4.800 2484.440 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2500.120 -4.800 2501.240 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2516.920 -4.800 2518.040 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2533.720 -4.800 2534.840 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 870.520 -4.800 871.640 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2550.520 -4.800 2551.640 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2567.320 -4.800 2568.440 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2584.120 -4.800 2585.240 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2600.920 -4.800 2602.040 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2617.720 -4.800 2618.840 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2634.520 -4.800 2635.640 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2651.320 -4.800 2652.440 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2668.120 -4.800 2669.240 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2684.920 -4.800 2686.040 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2701.720 -4.800 2702.840 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 887.320 -4.800 888.440 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2718.520 -4.800 2719.640 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2735.320 -4.800 2736.440 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2752.120 -4.800 2753.240 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2768.920 -4.800 2770.040 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2785.720 -4.800 2786.840 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2802.520 -4.800 2803.640 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2819.320 -4.800 2820.440 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2836.120 -4.800 2837.240 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 904.120 -4.800 905.240 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 920.920 -4.800 922.040 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 937.720 -4.800 938.840 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 954.520 -4.800 955.640 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 971.320 -4.800 972.440 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 988.120 -4.800 989.240 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1004.920 -4.800 1006.040 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1021.720 -4.800 1022.840 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 719.320 -4.800 720.440 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1038.520 -4.800 1039.640 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1055.320 -4.800 1056.440 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1072.120 -4.800 1073.240 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1088.920 -4.800 1090.040 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1105.720 -4.800 1106.840 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1122.520 -4.800 1123.640 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1139.320 -4.800 1140.440 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1156.120 -4.800 1157.240 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1172.920 -4.800 1174.040 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1189.720 -4.800 1190.840 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 736.120 -4.800 737.240 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1206.520 -4.800 1207.640 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1223.320 -4.800 1224.440 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1240.120 -4.800 1241.240 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1256.920 -4.800 1258.040 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1273.720 -4.800 1274.840 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1290.520 -4.800 1291.640 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1307.320 -4.800 1308.440 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1324.120 -4.800 1325.240 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1340.920 -4.800 1342.040 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1357.720 -4.800 1358.840 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 752.920 -4.800 754.040 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1374.520 -4.800 1375.640 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1391.320 -4.800 1392.440 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1408.120 -4.800 1409.240 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1424.920 -4.800 1426.040 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1441.720 -4.800 1442.840 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1458.520 -4.800 1459.640 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1475.320 -4.800 1476.440 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1492.120 -4.800 1493.240 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1508.920 -4.800 1510.040 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1525.720 -4.800 1526.840 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 769.720 -4.800 770.840 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1542.520 -4.800 1543.640 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1559.320 -4.800 1560.440 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1576.120 -4.800 1577.240 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1592.920 -4.800 1594.040 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1609.720 -4.800 1610.840 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1626.520 -4.800 1627.640 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1643.320 -4.800 1644.440 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1660.120 -4.800 1661.240 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1676.920 -4.800 1678.040 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1693.720 -4.800 1694.840 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 786.520 -4.800 787.640 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1710.520 -4.800 1711.640 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1727.320 -4.800 1728.440 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1744.120 -4.800 1745.240 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1760.920 -4.800 1762.040 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1777.720 -4.800 1778.840 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1794.520 -4.800 1795.640 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1811.320 -4.800 1812.440 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1828.120 -4.800 1829.240 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1844.920 -4.800 1846.040 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1861.720 -4.800 1862.840 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 803.320 -4.800 804.440 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1878.520 -4.800 1879.640 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1895.320 -4.800 1896.440 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1912.120 -4.800 1913.240 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1928.920 -4.800 1930.040 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1945.720 -4.800 1946.840 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1962.520 -4.800 1963.640 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1979.320 -4.800 1980.440 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1996.120 -4.800 1997.240 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2012.920 -4.800 2014.040 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2029.720 -4.800 2030.840 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 820.120 -4.800 821.240 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2046.520 -4.800 2047.640 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2063.320 -4.800 2064.440 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2080.120 -4.800 2081.240 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2096.920 -4.800 2098.040 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2113.720 -4.800 2114.840 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2130.520 -4.800 2131.640 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2147.320 -4.800 2148.440 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2164.120 -4.800 2165.240 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2180.920 -4.800 2182.040 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2197.720 -4.800 2198.840 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 836.920 -4.800 838.040 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2214.520 -4.800 2215.640 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2231.320 -4.800 2232.440 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2248.120 -4.800 2249.240 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2264.920 -4.800 2266.040 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2281.720 -4.800 2282.840 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2298.520 -4.800 2299.640 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2315.320 -4.800 2316.440 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2332.120 -4.800 2333.240 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2348.920 -4.800 2350.040 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2365.720 -4.800 2366.840 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 853.720 -4.800 854.840 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 708.120 -4.800 709.240 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2388.120 -4.800 2389.240 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2404.920 -4.800 2406.040 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2421.720 -4.800 2422.840 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2438.520 -4.800 2439.640 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2455.320 -4.800 2456.440 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2472.120 -4.800 2473.240 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2488.920 -4.800 2490.040 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2505.720 -4.800 2506.840 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2522.520 -4.800 2523.640 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2539.320 -4.800 2540.440 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 876.120 -4.800 877.240 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2556.120 -4.800 2557.240 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2572.920 -4.800 2574.040 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2589.720 -4.800 2590.840 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2606.520 -4.800 2607.640 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2623.320 -4.800 2624.440 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2640.120 -4.800 2641.240 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2656.920 -4.800 2658.040 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2673.720 -4.800 2674.840 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2690.520 -4.800 2691.640 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2707.320 -4.800 2708.440 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 892.920 -4.800 894.040 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2724.120 -4.800 2725.240 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2740.920 -4.800 2742.040 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2757.720 -4.800 2758.840 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2774.520 -4.800 2775.640 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2791.320 -4.800 2792.440 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2808.120 -4.800 2809.240 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2824.920 -4.800 2826.040 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2841.720 -4.800 2842.840 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 909.720 -4.800 910.840 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 926.520 -4.800 927.640 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 943.320 -4.800 944.440 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 960.120 -4.800 961.240 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 976.920 -4.800 978.040 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 993.720 -4.800 994.840 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1010.520 -4.800 1011.640 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1027.320 -4.800 1028.440 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 724.920 -4.800 726.040 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1044.120 -4.800 1045.240 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1060.920 -4.800 1062.040 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1077.720 -4.800 1078.840 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1094.520 -4.800 1095.640 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1111.320 -4.800 1112.440 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1128.120 -4.800 1129.240 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1144.920 -4.800 1146.040 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1161.720 -4.800 1162.840 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1178.520 -4.800 1179.640 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1195.320 -4.800 1196.440 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 741.720 -4.800 742.840 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1212.120 -4.800 1213.240 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1228.920 -4.800 1230.040 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1245.720 -4.800 1246.840 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1262.520 -4.800 1263.640 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1279.320 -4.800 1280.440 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1296.120 -4.800 1297.240 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1312.920 -4.800 1314.040 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1329.720 -4.800 1330.840 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1346.520 -4.800 1347.640 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1363.320 -4.800 1364.440 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 758.520 -4.800 759.640 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1380.120 -4.800 1381.240 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1396.920 -4.800 1398.040 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1413.720 -4.800 1414.840 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1430.520 -4.800 1431.640 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1447.320 -4.800 1448.440 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1464.120 -4.800 1465.240 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1480.920 -4.800 1482.040 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1497.720 -4.800 1498.840 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1514.520 -4.800 1515.640 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1531.320 -4.800 1532.440 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 775.320 -4.800 776.440 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1548.120 -4.800 1549.240 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1564.920 -4.800 1566.040 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1581.720 -4.800 1582.840 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1598.520 -4.800 1599.640 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1615.320 -4.800 1616.440 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1632.120 -4.800 1633.240 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1648.920 -4.800 1650.040 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1665.720 -4.800 1666.840 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1682.520 -4.800 1683.640 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1699.320 -4.800 1700.440 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 792.120 -4.800 793.240 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1716.120 -4.800 1717.240 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1732.920 -4.800 1734.040 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1749.720 -4.800 1750.840 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1766.520 -4.800 1767.640 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1783.320 -4.800 1784.440 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1800.120 -4.800 1801.240 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1816.920 -4.800 1818.040 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1833.720 -4.800 1834.840 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1850.520 -4.800 1851.640 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1867.320 -4.800 1868.440 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 808.920 -4.800 810.040 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1884.120 -4.800 1885.240 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1900.920 -4.800 1902.040 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1917.720 -4.800 1918.840 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1934.520 -4.800 1935.640 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1951.320 -4.800 1952.440 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1968.120 -4.800 1969.240 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1984.920 -4.800 1986.040 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2001.720 -4.800 2002.840 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2018.520 -4.800 2019.640 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2035.320 -4.800 2036.440 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 825.720 -4.800 826.840 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2052.120 -4.800 2053.240 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2068.920 -4.800 2070.040 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2085.720 -4.800 2086.840 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2102.520 -4.800 2103.640 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2119.320 -4.800 2120.440 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2136.120 -4.800 2137.240 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2152.920 -4.800 2154.040 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2169.720 -4.800 2170.840 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2186.520 -4.800 2187.640 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2203.320 -4.800 2204.440 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 842.520 -4.800 843.640 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2220.120 -4.800 2221.240 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2236.920 -4.800 2238.040 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2253.720 -4.800 2254.840 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2270.520 -4.800 2271.640 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2287.320 -4.800 2288.440 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2304.120 -4.800 2305.240 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2320.920 -4.800 2322.040 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2337.720 -4.800 2338.840 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2354.520 -4.800 2355.640 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2371.320 -4.800 2372.440 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 859.320 -4.800 860.440 2.400 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 713.720 -4.800 714.840 2.400 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2393.720 -4.800 2394.840 2.400 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2410.520 -4.800 2411.640 2.400 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2427.320 -4.800 2428.440 2.400 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2444.120 -4.800 2445.240 2.400 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2460.920 -4.800 2462.040 2.400 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2477.720 -4.800 2478.840 2.400 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2494.520 -4.800 2495.640 2.400 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2511.320 -4.800 2512.440 2.400 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2528.120 -4.800 2529.240 2.400 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2544.920 -4.800 2546.040 2.400 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 881.720 -4.800 882.840 2.400 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2561.720 -4.800 2562.840 2.400 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2578.520 -4.800 2579.640 2.400 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2595.320 -4.800 2596.440 2.400 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2612.120 -4.800 2613.240 2.400 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2628.920 -4.800 2630.040 2.400 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2645.720 -4.800 2646.840 2.400 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2662.520 -4.800 2663.640 2.400 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2679.320 -4.800 2680.440 2.400 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2696.120 -4.800 2697.240 2.400 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2712.920 -4.800 2714.040 2.400 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 898.520 -4.800 899.640 2.400 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2729.720 -4.800 2730.840 2.400 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2746.520 -4.800 2747.640 2.400 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2763.320 -4.800 2764.440 2.400 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2780.120 -4.800 2781.240 2.400 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2796.920 -4.800 2798.040 2.400 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2813.720 -4.800 2814.840 2.400 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2830.520 -4.800 2831.640 2.400 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2847.320 -4.800 2848.440 2.400 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 915.320 -4.800 916.440 2.400 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 932.120 -4.800 933.240 2.400 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 948.920 -4.800 950.040 2.400 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 965.720 -4.800 966.840 2.400 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 982.520 -4.800 983.640 2.400 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 999.320 -4.800 1000.440 2.400 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1016.120 -4.800 1017.240 2.400 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1032.920 -4.800 1034.040 2.400 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 730.520 -4.800 731.640 2.400 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1049.720 -4.800 1050.840 2.400 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1066.520 -4.800 1067.640 2.400 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1083.320 -4.800 1084.440 2.400 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1100.120 -4.800 1101.240 2.400 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1116.920 -4.800 1118.040 2.400 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1133.720 -4.800 1134.840 2.400 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1150.520 -4.800 1151.640 2.400 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1167.320 -4.800 1168.440 2.400 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1184.120 -4.800 1185.240 2.400 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1200.920 -4.800 1202.040 2.400 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 747.320 -4.800 748.440 2.400 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1217.720 -4.800 1218.840 2.400 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1234.520 -4.800 1235.640 2.400 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1251.320 -4.800 1252.440 2.400 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1268.120 -4.800 1269.240 2.400 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1284.920 -4.800 1286.040 2.400 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1301.720 -4.800 1302.840 2.400 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1318.520 -4.800 1319.640 2.400 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1335.320 -4.800 1336.440 2.400 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1352.120 -4.800 1353.240 2.400 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1368.920 -4.800 1370.040 2.400 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 764.120 -4.800 765.240 2.400 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1385.720 -4.800 1386.840 2.400 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1402.520 -4.800 1403.640 2.400 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1419.320 -4.800 1420.440 2.400 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1436.120 -4.800 1437.240 2.400 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1452.920 -4.800 1454.040 2.400 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1469.720 -4.800 1470.840 2.400 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1486.520 -4.800 1487.640 2.400 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1503.320 -4.800 1504.440 2.400 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1520.120 -4.800 1521.240 2.400 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1536.920 -4.800 1538.040 2.400 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 780.920 -4.800 782.040 2.400 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1553.720 -4.800 1554.840 2.400 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1570.520 -4.800 1571.640 2.400 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1587.320 -4.800 1588.440 2.400 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1604.120 -4.800 1605.240 2.400 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1620.920 -4.800 1622.040 2.400 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1637.720 -4.800 1638.840 2.400 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1654.520 -4.800 1655.640 2.400 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1671.320 -4.800 1672.440 2.400 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1688.120 -4.800 1689.240 2.400 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1704.920 -4.800 1706.040 2.400 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 797.720 -4.800 798.840 2.400 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1721.720 -4.800 1722.840 2.400 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1738.520 -4.800 1739.640 2.400 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1755.320 -4.800 1756.440 2.400 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1772.120 -4.800 1773.240 2.400 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1788.920 -4.800 1790.040 2.400 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1805.720 -4.800 1806.840 2.400 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1822.520 -4.800 1823.640 2.400 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1839.320 -4.800 1840.440 2.400 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1856.120 -4.800 1857.240 2.400 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1872.920 -4.800 1874.040 2.400 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 814.520 -4.800 815.640 2.400 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1889.720 -4.800 1890.840 2.400 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1906.520 -4.800 1907.640 2.400 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1923.320 -4.800 1924.440 2.400 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1940.120 -4.800 1941.240 2.400 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1956.920 -4.800 1958.040 2.400 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1973.720 -4.800 1974.840 2.400 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1990.520 -4.800 1991.640 2.400 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2007.320 -4.800 2008.440 2.400 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2024.120 -4.800 2025.240 2.400 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2040.920 -4.800 2042.040 2.400 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 831.320 -4.800 832.440 2.400 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2057.720 -4.800 2058.840 2.400 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2074.520 -4.800 2075.640 2.400 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2091.320 -4.800 2092.440 2.400 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2108.120 -4.800 2109.240 2.400 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2124.920 -4.800 2126.040 2.400 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2141.720 -4.800 2142.840 2.400 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2158.520 -4.800 2159.640 2.400 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2175.320 -4.800 2176.440 2.400 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2192.120 -4.800 2193.240 2.400 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2208.920 -4.800 2210.040 2.400 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 848.120 -4.800 849.240 2.400 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2225.720 -4.800 2226.840 2.400 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2242.520 -4.800 2243.640 2.400 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2259.320 -4.800 2260.440 2.400 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2276.120 -4.800 2277.240 2.400 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2292.920 -4.800 2294.040 2.400 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2309.720 -4.800 2310.840 2.400 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2326.520 -4.800 2327.640 2.400 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2343.320 -4.800 2344.440 2.400 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2360.120 -4.800 2361.240 2.400 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2376.920 -4.800 2378.040 2.400 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 864.920 -4.800 866.040 2.400 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2852.920 -4.800 2854.040 2.400 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2858.520 -4.800 2859.640 2.400 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2864.120 -4.800 2865.240 2.400 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2869.720 -4.800 2870.840 2.400 ;
    END
  END user_irq[2]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT -4.780 -3.420 -1.680 2986.540 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.780 -3.420 2985.100 -0.320 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.780 2983.440 2985.100 2986.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2982.000 -3.420 2985.100 2986.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 15.770 -8.220 18.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 105.770 -8.220 108.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 195.770 -8.220 198.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 285.770 -8.220 288.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 375.770 -8.220 378.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 465.770 -8.220 468.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 555.770 -8.220 558.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 645.770 -8.220 648.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 735.770 -8.220 738.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 825.770 -8.220 828.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 915.770 -8.220 918.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1005.770 -8.220 1008.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1095.770 -8.220 1098.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1185.770 -8.220 1188.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1275.770 -8.220 1278.870 1695.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1275.770 2284.660 1278.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1365.770 -8.220 1368.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1455.770 -8.220 1458.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1545.770 -8.220 1548.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1635.770 -8.220 1638.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1725.770 -8.220 1728.870 2247.650 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1725.770 2280.910 1728.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1815.770 -8.220 1818.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1905.770 -8.220 1908.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1995.770 -8.220 1998.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2085.770 -8.220 2088.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2175.770 -8.220 2178.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2265.770 -8.220 2268.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2355.770 -8.220 2358.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2445.770 -8.220 2448.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2535.770 -8.220 2538.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2625.770 -8.220 2628.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2715.770 -8.220 2718.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2805.770 -8.220 2808.870 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2895.770 -8.220 2898.870 2991.340 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 19.130 2989.900 22.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 109.130 2989.900 112.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 199.130 2989.900 202.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 289.130 2989.900 292.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 379.130 2989.900 382.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 469.130 2989.900 472.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 559.130 2989.900 562.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 649.130 2989.900 652.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 739.130 2989.900 742.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 829.130 2989.900 832.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 919.130 2989.900 922.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1009.130 2989.900 1012.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1099.130 2989.900 1102.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1189.130 2989.900 1192.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1279.130 2989.900 1282.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1369.130 2989.900 1372.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1459.130 2989.900 1462.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1549.130 2989.900 1552.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1639.130 2989.900 1642.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1729.130 2989.900 1732.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1819.130 2989.900 1822.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1909.130 2989.900 1912.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1999.130 2989.900 2002.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2089.130 2989.900 2092.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2179.130 2989.900 2182.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2269.130 2989.900 2272.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2359.130 2989.900 2362.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2449.130 2989.900 2452.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2539.130 2989.900 2542.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2629.130 2989.900 2632.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2719.130 2989.900 2722.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2809.130 2989.900 2812.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2899.130 2989.900 2902.230 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT -9.580 -8.220 -6.480 2991.340 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 -8.220 2989.900 -5.120 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2988.240 2989.900 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2986.800 -8.220 2989.900 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 34.370 -8.220 37.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 124.370 -8.220 127.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 214.370 -8.220 217.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 304.370 -8.220 307.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 394.370 -8.220 397.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 484.370 -8.220 487.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 574.370 -8.220 577.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 664.370 -8.220 667.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 754.370 -8.220 757.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 844.370 -8.220 847.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 934.370 -8.220 937.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1024.370 -8.220 1027.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1114.370 -8.220 1117.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1204.370 -8.220 1207.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1294.370 -8.220 1297.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1384.370 -8.220 1387.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1474.370 -8.220 1477.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1564.370 -8.220 1567.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1654.370 -8.220 1657.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1744.370 -8.220 1747.470 2247.650 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1744.370 2280.910 1747.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1834.370 -8.220 1837.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1924.370 -8.220 1927.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2014.370 -8.220 2017.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2104.370 -8.220 2107.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2194.370 -8.220 2197.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2284.370 -8.220 2287.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2374.370 -8.220 2377.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2464.370 -8.220 2467.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2554.370 -8.220 2557.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2644.370 -8.220 2647.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2734.370 -8.220 2737.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2824.370 -8.220 2827.470 2991.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2914.370 -8.220 2917.470 2991.340 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 49.130 2989.900 52.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 139.130 2989.900 142.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 229.130 2989.900 232.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 319.130 2989.900 322.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 409.130 2989.900 412.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 499.130 2989.900 502.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 589.130 2989.900 592.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 679.130 2989.900 682.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 769.130 2989.900 772.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 859.130 2989.900 862.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 949.130 2989.900 952.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1039.130 2989.900 1042.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1129.130 2989.900 1132.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1219.130 2989.900 1222.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1309.130 2989.900 1312.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1399.130 2989.900 1402.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1489.130 2989.900 1492.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1579.130 2989.900 1582.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1669.130 2989.900 1672.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1759.130 2989.900 1762.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1849.130 2989.900 1852.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 1939.130 2989.900 1942.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2029.130 2989.900 2032.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2119.130 2989.900 2122.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2209.130 2989.900 2212.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2299.130 2989.900 2302.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2389.130 2989.900 2392.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2479.130 2989.900 2482.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2569.130 2989.900 2572.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2659.130 2989.900 2662.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2749.130 2989.900 2752.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2839.130 2989.900 2842.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -9.580 2929.130 2989.900 2932.230 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 108.920 -4.800 110.040 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 114.520 -4.800 115.640 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 120.120 -4.800 121.240 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 142.520 -4.800 143.640 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 332.920 -4.800 334.040 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 349.720 -4.800 350.840 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 366.520 -4.800 367.640 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 383.320 -4.800 384.440 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 400.120 -4.800 401.240 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 416.920 -4.800 418.040 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 433.720 -4.800 434.840 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 450.520 -4.800 451.640 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 467.320 -4.800 468.440 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 484.120 -4.800 485.240 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 164.920 -4.800 166.040 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 500.920 -4.800 502.040 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 517.720 -4.800 518.840 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 534.520 -4.800 535.640 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 551.320 -4.800 552.440 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 568.120 -4.800 569.240 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 584.920 -4.800 586.040 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 601.720 -4.800 602.840 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 618.520 -4.800 619.640 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 635.320 -4.800 636.440 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 652.120 -4.800 653.240 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 187.320 -4.800 188.440 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 668.920 -4.800 670.040 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 685.720 -4.800 686.840 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 209.720 -4.800 210.840 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 232.120 -4.800 233.240 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 248.920 -4.800 250.040 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 265.720 -4.800 266.840 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 282.520 -4.800 283.640 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 299.320 -4.800 300.440 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 316.120 -4.800 317.240 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 125.720 -4.800 126.840 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 148.120 -4.800 149.240 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 338.520 -4.800 339.640 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 355.320 -4.800 356.440 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 372.120 -4.800 373.240 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 388.920 -4.800 390.040 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 405.720 -4.800 406.840 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 422.520 -4.800 423.640 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 439.320 -4.800 440.440 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 456.120 -4.800 457.240 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 472.920 -4.800 474.040 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 489.720 -4.800 490.840 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 170.520 -4.800 171.640 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 506.520 -4.800 507.640 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 523.320 -4.800 524.440 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 540.120 -4.800 541.240 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 556.920 -4.800 558.040 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 573.720 -4.800 574.840 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 590.520 -4.800 591.640 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 607.320 -4.800 608.440 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 624.120 -4.800 625.240 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 640.920 -4.800 642.040 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 657.720 -4.800 658.840 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 192.920 -4.800 194.040 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 674.520 -4.800 675.640 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 691.320 -4.800 692.440 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 215.320 -4.800 216.440 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 237.720 -4.800 238.840 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 254.520 -4.800 255.640 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 271.320 -4.800 272.440 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 288.120 -4.800 289.240 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 304.920 -4.800 306.040 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 321.720 -4.800 322.840 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 153.720 -4.800 154.840 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 344.120 -4.800 345.240 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 360.920 -4.800 362.040 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 377.720 -4.800 378.840 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 394.520 -4.800 395.640 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 411.320 -4.800 412.440 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 428.120 -4.800 429.240 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 444.920 -4.800 446.040 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 461.720 -4.800 462.840 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 478.520 -4.800 479.640 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 495.320 -4.800 496.440 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 176.120 -4.800 177.240 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 512.120 -4.800 513.240 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 528.920 -4.800 530.040 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 545.720 -4.800 546.840 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 562.520 -4.800 563.640 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 579.320 -4.800 580.440 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 596.120 -4.800 597.240 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 612.920 -4.800 614.040 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 629.720 -4.800 630.840 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 646.520 -4.800 647.640 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 663.320 -4.800 664.440 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 198.520 -4.800 199.640 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 680.120 -4.800 681.240 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 696.920 -4.800 698.040 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 220.920 -4.800 222.040 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 243.320 -4.800 244.440 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 260.120 -4.800 261.240 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 276.920 -4.800 278.040 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 293.720 -4.800 294.840 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 310.520 -4.800 311.640 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 327.320 -4.800 328.440 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 159.320 -4.800 160.440 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 181.720 -4.800 182.840 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 204.120 -4.800 205.240 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 226.520 -4.800 227.640 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 131.320 -4.800 132.440 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 136.920 -4.800 138.040 2.400 ;
    END
  END wbs_we_i
  OBS
      LAYER Metal1 ;
        RECT 344.490 46.070 2785.910 2286.890 ;
      LAYER Metal2 ;
        RECT 12.460 2977.500 48.700 2978.500 ;
        RECT 50.420 2977.500 131.020 2978.500 ;
        RECT 132.740 2977.500 213.340 2978.500 ;
        RECT 215.060 2977.500 295.660 2978.500 ;
        RECT 297.380 2977.500 377.980 2978.500 ;
        RECT 379.700 2977.500 460.300 2978.500 ;
        RECT 462.020 2977.500 542.620 2978.500 ;
        RECT 544.340 2977.500 624.940 2978.500 ;
        RECT 626.660 2977.500 707.260 2978.500 ;
        RECT 708.980 2977.500 789.580 2978.500 ;
        RECT 791.300 2977.500 871.900 2978.500 ;
        RECT 873.620 2977.500 954.220 2978.500 ;
        RECT 955.940 2977.500 1036.540 2978.500 ;
        RECT 1038.260 2977.500 1118.860 2978.500 ;
        RECT 1120.580 2977.500 1201.180 2978.500 ;
        RECT 1202.900 2977.500 1283.500 2978.500 ;
        RECT 1285.220 2977.500 1365.820 2978.500 ;
        RECT 1367.540 2977.500 1448.140 2978.500 ;
        RECT 1449.860 2977.500 1530.460 2978.500 ;
        RECT 1532.180 2977.500 1612.780 2978.500 ;
        RECT 1614.500 2977.500 1695.100 2978.500 ;
        RECT 1696.820 2977.500 1777.420 2978.500 ;
        RECT 1779.140 2977.500 1859.740 2978.500 ;
        RECT 1861.460 2977.500 1942.060 2978.500 ;
        RECT 1943.780 2977.500 2024.380 2978.500 ;
        RECT 2026.100 2977.500 2106.700 2978.500 ;
        RECT 2108.420 2977.500 2189.020 2978.500 ;
        RECT 2190.740 2977.500 2271.340 2978.500 ;
        RECT 2273.060 2977.500 2353.660 2978.500 ;
        RECT 2355.380 2977.500 2435.980 2978.500 ;
        RECT 2437.700 2977.500 2518.300 2978.500 ;
        RECT 2520.020 2977.500 2600.620 2978.500 ;
        RECT 2602.340 2977.500 2682.940 2978.500 ;
        RECT 2684.660 2977.500 2765.260 2978.500 ;
        RECT 2766.980 2977.500 2847.580 2978.500 ;
        RECT 2849.300 2977.500 2929.900 2978.500 ;
        RECT 2931.620 2977.500 2970.100 2978.500 ;
        RECT 12.460 2.700 2970.100 2977.500 ;
        RECT 12.460 1.820 108.620 2.700 ;
        RECT 110.340 1.820 114.220 2.700 ;
        RECT 115.940 1.820 119.820 2.700 ;
        RECT 121.540 1.820 125.420 2.700 ;
        RECT 127.140 1.820 131.020 2.700 ;
        RECT 132.740 1.820 136.620 2.700 ;
        RECT 138.340 1.820 142.220 2.700 ;
        RECT 143.940 1.820 147.820 2.700 ;
        RECT 149.540 1.820 153.420 2.700 ;
        RECT 155.140 1.820 159.020 2.700 ;
        RECT 160.740 1.820 164.620 2.700 ;
        RECT 166.340 1.820 170.220 2.700 ;
        RECT 171.940 1.820 175.820 2.700 ;
        RECT 177.540 1.820 181.420 2.700 ;
        RECT 183.140 1.820 187.020 2.700 ;
        RECT 188.740 1.820 192.620 2.700 ;
        RECT 194.340 1.820 198.220 2.700 ;
        RECT 199.940 1.820 203.820 2.700 ;
        RECT 205.540 1.820 209.420 2.700 ;
        RECT 211.140 1.820 215.020 2.700 ;
        RECT 216.740 1.820 220.620 2.700 ;
        RECT 222.340 1.820 226.220 2.700 ;
        RECT 227.940 1.820 231.820 2.700 ;
        RECT 233.540 1.820 237.420 2.700 ;
        RECT 239.140 1.820 243.020 2.700 ;
        RECT 244.740 1.820 248.620 2.700 ;
        RECT 250.340 1.820 254.220 2.700 ;
        RECT 255.940 1.820 259.820 2.700 ;
        RECT 261.540 1.820 265.420 2.700 ;
        RECT 267.140 1.820 271.020 2.700 ;
        RECT 272.740 1.820 276.620 2.700 ;
        RECT 278.340 1.820 282.220 2.700 ;
        RECT 283.940 1.820 287.820 2.700 ;
        RECT 289.540 1.820 293.420 2.700 ;
        RECT 295.140 1.820 299.020 2.700 ;
        RECT 300.740 1.820 304.620 2.700 ;
        RECT 306.340 1.820 310.220 2.700 ;
        RECT 311.940 1.820 315.820 2.700 ;
        RECT 317.540 1.820 321.420 2.700 ;
        RECT 323.140 1.820 327.020 2.700 ;
        RECT 328.740 1.820 332.620 2.700 ;
        RECT 334.340 1.820 338.220 2.700 ;
        RECT 339.940 1.820 343.820 2.700 ;
        RECT 345.540 1.820 349.420 2.700 ;
        RECT 351.140 1.820 355.020 2.700 ;
        RECT 356.740 1.820 360.620 2.700 ;
        RECT 362.340 1.820 366.220 2.700 ;
        RECT 367.940 1.820 371.820 2.700 ;
        RECT 373.540 1.820 377.420 2.700 ;
        RECT 379.140 1.820 383.020 2.700 ;
        RECT 384.740 1.820 388.620 2.700 ;
        RECT 390.340 1.820 394.220 2.700 ;
        RECT 395.940 1.820 399.820 2.700 ;
        RECT 401.540 1.820 405.420 2.700 ;
        RECT 407.140 1.820 411.020 2.700 ;
        RECT 412.740 1.820 416.620 2.700 ;
        RECT 418.340 1.820 422.220 2.700 ;
        RECT 423.940 1.820 427.820 2.700 ;
        RECT 429.540 1.820 433.420 2.700 ;
        RECT 435.140 1.820 439.020 2.700 ;
        RECT 440.740 1.820 444.620 2.700 ;
        RECT 446.340 1.820 450.220 2.700 ;
        RECT 451.940 1.820 455.820 2.700 ;
        RECT 457.540 1.820 461.420 2.700 ;
        RECT 463.140 1.820 467.020 2.700 ;
        RECT 468.740 1.820 472.620 2.700 ;
        RECT 474.340 1.820 478.220 2.700 ;
        RECT 479.940 1.820 483.820 2.700 ;
        RECT 485.540 1.820 489.420 2.700 ;
        RECT 491.140 1.820 495.020 2.700 ;
        RECT 496.740 1.820 500.620 2.700 ;
        RECT 502.340 1.820 506.220 2.700 ;
        RECT 507.940 1.820 511.820 2.700 ;
        RECT 513.540 1.820 517.420 2.700 ;
        RECT 519.140 1.820 523.020 2.700 ;
        RECT 524.740 1.820 528.620 2.700 ;
        RECT 530.340 1.820 534.220 2.700 ;
        RECT 535.940 1.820 539.820 2.700 ;
        RECT 541.540 1.820 545.420 2.700 ;
        RECT 547.140 1.820 551.020 2.700 ;
        RECT 552.740 1.820 556.620 2.700 ;
        RECT 558.340 1.820 562.220 2.700 ;
        RECT 563.940 1.820 567.820 2.700 ;
        RECT 569.540 1.820 573.420 2.700 ;
        RECT 575.140 1.820 579.020 2.700 ;
        RECT 580.740 1.820 584.620 2.700 ;
        RECT 586.340 1.820 590.220 2.700 ;
        RECT 591.940 1.820 595.820 2.700 ;
        RECT 597.540 1.820 601.420 2.700 ;
        RECT 603.140 1.820 607.020 2.700 ;
        RECT 608.740 1.820 612.620 2.700 ;
        RECT 614.340 1.820 618.220 2.700 ;
        RECT 619.940 1.820 623.820 2.700 ;
        RECT 625.540 1.820 629.420 2.700 ;
        RECT 631.140 1.820 635.020 2.700 ;
        RECT 636.740 1.820 640.620 2.700 ;
        RECT 642.340 1.820 646.220 2.700 ;
        RECT 647.940 1.820 651.820 2.700 ;
        RECT 653.540 1.820 657.420 2.700 ;
        RECT 659.140 1.820 663.020 2.700 ;
        RECT 664.740 1.820 668.620 2.700 ;
        RECT 670.340 1.820 674.220 2.700 ;
        RECT 675.940 1.820 679.820 2.700 ;
        RECT 681.540 1.820 685.420 2.700 ;
        RECT 687.140 1.820 691.020 2.700 ;
        RECT 692.740 1.820 696.620 2.700 ;
        RECT 698.340 1.820 702.220 2.700 ;
        RECT 703.940 1.820 707.820 2.700 ;
        RECT 709.540 1.820 713.420 2.700 ;
        RECT 715.140 1.820 719.020 2.700 ;
        RECT 720.740 1.820 724.620 2.700 ;
        RECT 726.340 1.820 730.220 2.700 ;
        RECT 731.940 1.820 735.820 2.700 ;
        RECT 737.540 1.820 741.420 2.700 ;
        RECT 743.140 1.820 747.020 2.700 ;
        RECT 748.740 1.820 752.620 2.700 ;
        RECT 754.340 1.820 758.220 2.700 ;
        RECT 759.940 1.820 763.820 2.700 ;
        RECT 765.540 1.820 769.420 2.700 ;
        RECT 771.140 1.820 775.020 2.700 ;
        RECT 776.740 1.820 780.620 2.700 ;
        RECT 782.340 1.820 786.220 2.700 ;
        RECT 787.940 1.820 791.820 2.700 ;
        RECT 793.540 1.820 797.420 2.700 ;
        RECT 799.140 1.820 803.020 2.700 ;
        RECT 804.740 1.820 808.620 2.700 ;
        RECT 810.340 1.820 814.220 2.700 ;
        RECT 815.940 1.820 819.820 2.700 ;
        RECT 821.540 1.820 825.420 2.700 ;
        RECT 827.140 1.820 831.020 2.700 ;
        RECT 832.740 1.820 836.620 2.700 ;
        RECT 838.340 1.820 842.220 2.700 ;
        RECT 843.940 1.820 847.820 2.700 ;
        RECT 849.540 1.820 853.420 2.700 ;
        RECT 855.140 1.820 859.020 2.700 ;
        RECT 860.740 1.820 864.620 2.700 ;
        RECT 866.340 1.820 870.220 2.700 ;
        RECT 871.940 1.820 875.820 2.700 ;
        RECT 877.540 1.820 881.420 2.700 ;
        RECT 883.140 1.820 887.020 2.700 ;
        RECT 888.740 1.820 892.620 2.700 ;
        RECT 894.340 1.820 898.220 2.700 ;
        RECT 899.940 1.820 903.820 2.700 ;
        RECT 905.540 1.820 909.420 2.700 ;
        RECT 911.140 1.820 915.020 2.700 ;
        RECT 916.740 1.820 920.620 2.700 ;
        RECT 922.340 1.820 926.220 2.700 ;
        RECT 927.940 1.820 931.820 2.700 ;
        RECT 933.540 1.820 937.420 2.700 ;
        RECT 939.140 1.820 943.020 2.700 ;
        RECT 944.740 1.820 948.620 2.700 ;
        RECT 950.340 1.820 954.220 2.700 ;
        RECT 955.940 1.820 959.820 2.700 ;
        RECT 961.540 1.820 965.420 2.700 ;
        RECT 967.140 1.820 971.020 2.700 ;
        RECT 972.740 1.820 976.620 2.700 ;
        RECT 978.340 1.820 982.220 2.700 ;
        RECT 983.940 1.820 987.820 2.700 ;
        RECT 989.540 1.820 993.420 2.700 ;
        RECT 995.140 1.820 999.020 2.700 ;
        RECT 1000.740 1.820 1004.620 2.700 ;
        RECT 1006.340 1.820 1010.220 2.700 ;
        RECT 1011.940 1.820 1015.820 2.700 ;
        RECT 1017.540 1.820 1021.420 2.700 ;
        RECT 1023.140 1.820 1027.020 2.700 ;
        RECT 1028.740 1.820 1032.620 2.700 ;
        RECT 1034.340 1.820 1038.220 2.700 ;
        RECT 1039.940 1.820 1043.820 2.700 ;
        RECT 1045.540 1.820 1049.420 2.700 ;
        RECT 1051.140 1.820 1055.020 2.700 ;
        RECT 1056.740 1.820 1060.620 2.700 ;
        RECT 1062.340 1.820 1066.220 2.700 ;
        RECT 1067.940 1.820 1071.820 2.700 ;
        RECT 1073.540 1.820 1077.420 2.700 ;
        RECT 1079.140 1.820 1083.020 2.700 ;
        RECT 1084.740 1.820 1088.620 2.700 ;
        RECT 1090.340 1.820 1094.220 2.700 ;
        RECT 1095.940 1.820 1099.820 2.700 ;
        RECT 1101.540 1.820 1105.420 2.700 ;
        RECT 1107.140 1.820 1111.020 2.700 ;
        RECT 1112.740 1.820 1116.620 2.700 ;
        RECT 1118.340 1.820 1122.220 2.700 ;
        RECT 1123.940 1.820 1127.820 2.700 ;
        RECT 1129.540 1.820 1133.420 2.700 ;
        RECT 1135.140 1.820 1139.020 2.700 ;
        RECT 1140.740 1.820 1144.620 2.700 ;
        RECT 1146.340 1.820 1150.220 2.700 ;
        RECT 1151.940 1.820 1155.820 2.700 ;
        RECT 1157.540 1.820 1161.420 2.700 ;
        RECT 1163.140 1.820 1167.020 2.700 ;
        RECT 1168.740 1.820 1172.620 2.700 ;
        RECT 1174.340 1.820 1178.220 2.700 ;
        RECT 1179.940 1.820 1183.820 2.700 ;
        RECT 1185.540 1.820 1189.420 2.700 ;
        RECT 1191.140 1.820 1195.020 2.700 ;
        RECT 1196.740 1.820 1200.620 2.700 ;
        RECT 1202.340 1.820 1206.220 2.700 ;
        RECT 1207.940 1.820 1211.820 2.700 ;
        RECT 1213.540 1.820 1217.420 2.700 ;
        RECT 1219.140 1.820 1223.020 2.700 ;
        RECT 1224.740 1.820 1228.620 2.700 ;
        RECT 1230.340 1.820 1234.220 2.700 ;
        RECT 1235.940 1.820 1239.820 2.700 ;
        RECT 1241.540 1.820 1245.420 2.700 ;
        RECT 1247.140 1.820 1251.020 2.700 ;
        RECT 1252.740 1.820 1256.620 2.700 ;
        RECT 1258.340 1.820 1262.220 2.700 ;
        RECT 1263.940 1.820 1267.820 2.700 ;
        RECT 1269.540 1.820 1273.420 2.700 ;
        RECT 1275.140 1.820 1279.020 2.700 ;
        RECT 1280.740 1.820 1284.620 2.700 ;
        RECT 1286.340 1.820 1290.220 2.700 ;
        RECT 1291.940 1.820 1295.820 2.700 ;
        RECT 1297.540 1.820 1301.420 2.700 ;
        RECT 1303.140 1.820 1307.020 2.700 ;
        RECT 1308.740 1.820 1312.620 2.700 ;
        RECT 1314.340 1.820 1318.220 2.700 ;
        RECT 1319.940 1.820 1323.820 2.700 ;
        RECT 1325.540 1.820 1329.420 2.700 ;
        RECT 1331.140 1.820 1335.020 2.700 ;
        RECT 1336.740 1.820 1340.620 2.700 ;
        RECT 1342.340 1.820 1346.220 2.700 ;
        RECT 1347.940 1.820 1351.820 2.700 ;
        RECT 1353.540 1.820 1357.420 2.700 ;
        RECT 1359.140 1.820 1363.020 2.700 ;
        RECT 1364.740 1.820 1368.620 2.700 ;
        RECT 1370.340 1.820 1374.220 2.700 ;
        RECT 1375.940 1.820 1379.820 2.700 ;
        RECT 1381.540 1.820 1385.420 2.700 ;
        RECT 1387.140 1.820 1391.020 2.700 ;
        RECT 1392.740 1.820 1396.620 2.700 ;
        RECT 1398.340 1.820 1402.220 2.700 ;
        RECT 1403.940 1.820 1407.820 2.700 ;
        RECT 1409.540 1.820 1413.420 2.700 ;
        RECT 1415.140 1.820 1419.020 2.700 ;
        RECT 1420.740 1.820 1424.620 2.700 ;
        RECT 1426.340 1.820 1430.220 2.700 ;
        RECT 1431.940 1.820 1435.820 2.700 ;
        RECT 1437.540 1.820 1441.420 2.700 ;
        RECT 1443.140 1.820 1447.020 2.700 ;
        RECT 1448.740 1.820 1452.620 2.700 ;
        RECT 1454.340 1.820 1458.220 2.700 ;
        RECT 1459.940 1.820 1463.820 2.700 ;
        RECT 1465.540 1.820 1469.420 2.700 ;
        RECT 1471.140 1.820 1475.020 2.700 ;
        RECT 1476.740 1.820 1480.620 2.700 ;
        RECT 1482.340 1.820 1486.220 2.700 ;
        RECT 1487.940 1.820 1491.820 2.700 ;
        RECT 1493.540 1.820 1497.420 2.700 ;
        RECT 1499.140 1.820 1503.020 2.700 ;
        RECT 1504.740 1.820 1508.620 2.700 ;
        RECT 1510.340 1.820 1514.220 2.700 ;
        RECT 1515.940 1.820 1519.820 2.700 ;
        RECT 1521.540 1.820 1525.420 2.700 ;
        RECT 1527.140 1.820 1531.020 2.700 ;
        RECT 1532.740 1.820 1536.620 2.700 ;
        RECT 1538.340 1.820 1542.220 2.700 ;
        RECT 1543.940 1.820 1547.820 2.700 ;
        RECT 1549.540 1.820 1553.420 2.700 ;
        RECT 1555.140 1.820 1559.020 2.700 ;
        RECT 1560.740 1.820 1564.620 2.700 ;
        RECT 1566.340 1.820 1570.220 2.700 ;
        RECT 1571.940 1.820 1575.820 2.700 ;
        RECT 1577.540 1.820 1581.420 2.700 ;
        RECT 1583.140 1.820 1587.020 2.700 ;
        RECT 1588.740 1.820 1592.620 2.700 ;
        RECT 1594.340 1.820 1598.220 2.700 ;
        RECT 1599.940 1.820 1603.820 2.700 ;
        RECT 1605.540 1.820 1609.420 2.700 ;
        RECT 1611.140 1.820 1615.020 2.700 ;
        RECT 1616.740 1.820 1620.620 2.700 ;
        RECT 1622.340 1.820 1626.220 2.700 ;
        RECT 1627.940 1.820 1631.820 2.700 ;
        RECT 1633.540 1.820 1637.420 2.700 ;
        RECT 1639.140 1.820 1643.020 2.700 ;
        RECT 1644.740 1.820 1648.620 2.700 ;
        RECT 1650.340 1.820 1654.220 2.700 ;
        RECT 1655.940 1.820 1659.820 2.700 ;
        RECT 1661.540 1.820 1665.420 2.700 ;
        RECT 1667.140 1.820 1671.020 2.700 ;
        RECT 1672.740 1.820 1676.620 2.700 ;
        RECT 1678.340 1.820 1682.220 2.700 ;
        RECT 1683.940 1.820 1687.820 2.700 ;
        RECT 1689.540 1.820 1693.420 2.700 ;
        RECT 1695.140 1.820 1699.020 2.700 ;
        RECT 1700.740 1.820 1704.620 2.700 ;
        RECT 1706.340 1.820 1710.220 2.700 ;
        RECT 1711.940 1.820 1715.820 2.700 ;
        RECT 1717.540 1.820 1721.420 2.700 ;
        RECT 1723.140 1.820 1727.020 2.700 ;
        RECT 1728.740 1.820 1732.620 2.700 ;
        RECT 1734.340 1.820 1738.220 2.700 ;
        RECT 1739.940 1.820 1743.820 2.700 ;
        RECT 1745.540 1.820 1749.420 2.700 ;
        RECT 1751.140 1.820 1755.020 2.700 ;
        RECT 1756.740 1.820 1760.620 2.700 ;
        RECT 1762.340 1.820 1766.220 2.700 ;
        RECT 1767.940 1.820 1771.820 2.700 ;
        RECT 1773.540 1.820 1777.420 2.700 ;
        RECT 1779.140 1.820 1783.020 2.700 ;
        RECT 1784.740 1.820 1788.620 2.700 ;
        RECT 1790.340 1.820 1794.220 2.700 ;
        RECT 1795.940 1.820 1799.820 2.700 ;
        RECT 1801.540 1.820 1805.420 2.700 ;
        RECT 1807.140 1.820 1811.020 2.700 ;
        RECT 1812.740 1.820 1816.620 2.700 ;
        RECT 1818.340 1.820 1822.220 2.700 ;
        RECT 1823.940 1.820 1827.820 2.700 ;
        RECT 1829.540 1.820 1833.420 2.700 ;
        RECT 1835.140 1.820 1839.020 2.700 ;
        RECT 1840.740 1.820 1844.620 2.700 ;
        RECT 1846.340 1.820 1850.220 2.700 ;
        RECT 1851.940 1.820 1855.820 2.700 ;
        RECT 1857.540 1.820 1861.420 2.700 ;
        RECT 1863.140 1.820 1867.020 2.700 ;
        RECT 1868.740 1.820 1872.620 2.700 ;
        RECT 1874.340 1.820 1878.220 2.700 ;
        RECT 1879.940 1.820 1883.820 2.700 ;
        RECT 1885.540 1.820 1889.420 2.700 ;
        RECT 1891.140 1.820 1895.020 2.700 ;
        RECT 1896.740 1.820 1900.620 2.700 ;
        RECT 1902.340 1.820 1906.220 2.700 ;
        RECT 1907.940 1.820 1911.820 2.700 ;
        RECT 1913.540 1.820 1917.420 2.700 ;
        RECT 1919.140 1.820 1923.020 2.700 ;
        RECT 1924.740 1.820 1928.620 2.700 ;
        RECT 1930.340 1.820 1934.220 2.700 ;
        RECT 1935.940 1.820 1939.820 2.700 ;
        RECT 1941.540 1.820 1945.420 2.700 ;
        RECT 1947.140 1.820 1951.020 2.700 ;
        RECT 1952.740 1.820 1956.620 2.700 ;
        RECT 1958.340 1.820 1962.220 2.700 ;
        RECT 1963.940 1.820 1967.820 2.700 ;
        RECT 1969.540 1.820 1973.420 2.700 ;
        RECT 1975.140 1.820 1979.020 2.700 ;
        RECT 1980.740 1.820 1984.620 2.700 ;
        RECT 1986.340 1.820 1990.220 2.700 ;
        RECT 1991.940 1.820 1995.820 2.700 ;
        RECT 1997.540 1.820 2001.420 2.700 ;
        RECT 2003.140 1.820 2007.020 2.700 ;
        RECT 2008.740 1.820 2012.620 2.700 ;
        RECT 2014.340 1.820 2018.220 2.700 ;
        RECT 2019.940 1.820 2023.820 2.700 ;
        RECT 2025.540 1.820 2029.420 2.700 ;
        RECT 2031.140 1.820 2035.020 2.700 ;
        RECT 2036.740 1.820 2040.620 2.700 ;
        RECT 2042.340 1.820 2046.220 2.700 ;
        RECT 2047.940 1.820 2051.820 2.700 ;
        RECT 2053.540 1.820 2057.420 2.700 ;
        RECT 2059.140 1.820 2063.020 2.700 ;
        RECT 2064.740 1.820 2068.620 2.700 ;
        RECT 2070.340 1.820 2074.220 2.700 ;
        RECT 2075.940 1.820 2079.820 2.700 ;
        RECT 2081.540 1.820 2085.420 2.700 ;
        RECT 2087.140 1.820 2091.020 2.700 ;
        RECT 2092.740 1.820 2096.620 2.700 ;
        RECT 2098.340 1.820 2102.220 2.700 ;
        RECT 2103.940 1.820 2107.820 2.700 ;
        RECT 2109.540 1.820 2113.420 2.700 ;
        RECT 2115.140 1.820 2119.020 2.700 ;
        RECT 2120.740 1.820 2124.620 2.700 ;
        RECT 2126.340 1.820 2130.220 2.700 ;
        RECT 2131.940 1.820 2135.820 2.700 ;
        RECT 2137.540 1.820 2141.420 2.700 ;
        RECT 2143.140 1.820 2147.020 2.700 ;
        RECT 2148.740 1.820 2152.620 2.700 ;
        RECT 2154.340 1.820 2158.220 2.700 ;
        RECT 2159.940 1.820 2163.820 2.700 ;
        RECT 2165.540 1.820 2169.420 2.700 ;
        RECT 2171.140 1.820 2175.020 2.700 ;
        RECT 2176.740 1.820 2180.620 2.700 ;
        RECT 2182.340 1.820 2186.220 2.700 ;
        RECT 2187.940 1.820 2191.820 2.700 ;
        RECT 2193.540 1.820 2197.420 2.700 ;
        RECT 2199.140 1.820 2203.020 2.700 ;
        RECT 2204.740 1.820 2208.620 2.700 ;
        RECT 2210.340 1.820 2214.220 2.700 ;
        RECT 2215.940 1.820 2219.820 2.700 ;
        RECT 2221.540 1.820 2225.420 2.700 ;
        RECT 2227.140 1.820 2231.020 2.700 ;
        RECT 2232.740 1.820 2236.620 2.700 ;
        RECT 2238.340 1.820 2242.220 2.700 ;
        RECT 2243.940 1.820 2247.820 2.700 ;
        RECT 2249.540 1.820 2253.420 2.700 ;
        RECT 2255.140 1.820 2259.020 2.700 ;
        RECT 2260.740 1.820 2264.620 2.700 ;
        RECT 2266.340 1.820 2270.220 2.700 ;
        RECT 2271.940 1.820 2275.820 2.700 ;
        RECT 2277.540 1.820 2281.420 2.700 ;
        RECT 2283.140 1.820 2287.020 2.700 ;
        RECT 2288.740 1.820 2292.620 2.700 ;
        RECT 2294.340 1.820 2298.220 2.700 ;
        RECT 2299.940 1.820 2303.820 2.700 ;
        RECT 2305.540 1.820 2309.420 2.700 ;
        RECT 2311.140 1.820 2315.020 2.700 ;
        RECT 2316.740 1.820 2320.620 2.700 ;
        RECT 2322.340 1.820 2326.220 2.700 ;
        RECT 2327.940 1.820 2331.820 2.700 ;
        RECT 2333.540 1.820 2337.420 2.700 ;
        RECT 2339.140 1.820 2343.020 2.700 ;
        RECT 2344.740 1.820 2348.620 2.700 ;
        RECT 2350.340 1.820 2354.220 2.700 ;
        RECT 2355.940 1.820 2359.820 2.700 ;
        RECT 2361.540 1.820 2365.420 2.700 ;
        RECT 2367.140 1.820 2371.020 2.700 ;
        RECT 2372.740 1.820 2376.620 2.700 ;
        RECT 2378.340 1.820 2382.220 2.700 ;
        RECT 2383.940 1.820 2387.820 2.700 ;
        RECT 2389.540 1.820 2393.420 2.700 ;
        RECT 2395.140 1.820 2399.020 2.700 ;
        RECT 2400.740 1.820 2404.620 2.700 ;
        RECT 2406.340 1.820 2410.220 2.700 ;
        RECT 2411.940 1.820 2415.820 2.700 ;
        RECT 2417.540 1.820 2421.420 2.700 ;
        RECT 2423.140 1.820 2427.020 2.700 ;
        RECT 2428.740 1.820 2432.620 2.700 ;
        RECT 2434.340 1.820 2438.220 2.700 ;
        RECT 2439.940 1.820 2443.820 2.700 ;
        RECT 2445.540 1.820 2449.420 2.700 ;
        RECT 2451.140 1.820 2455.020 2.700 ;
        RECT 2456.740 1.820 2460.620 2.700 ;
        RECT 2462.340 1.820 2466.220 2.700 ;
        RECT 2467.940 1.820 2471.820 2.700 ;
        RECT 2473.540 1.820 2477.420 2.700 ;
        RECT 2479.140 1.820 2483.020 2.700 ;
        RECT 2484.740 1.820 2488.620 2.700 ;
        RECT 2490.340 1.820 2494.220 2.700 ;
        RECT 2495.940 1.820 2499.820 2.700 ;
        RECT 2501.540 1.820 2505.420 2.700 ;
        RECT 2507.140 1.820 2511.020 2.700 ;
        RECT 2512.740 1.820 2516.620 2.700 ;
        RECT 2518.340 1.820 2522.220 2.700 ;
        RECT 2523.940 1.820 2527.820 2.700 ;
        RECT 2529.540 1.820 2533.420 2.700 ;
        RECT 2535.140 1.820 2539.020 2.700 ;
        RECT 2540.740 1.820 2544.620 2.700 ;
        RECT 2546.340 1.820 2550.220 2.700 ;
        RECT 2551.940 1.820 2555.820 2.700 ;
        RECT 2557.540 1.820 2561.420 2.700 ;
        RECT 2563.140 1.820 2567.020 2.700 ;
        RECT 2568.740 1.820 2572.620 2.700 ;
        RECT 2574.340 1.820 2578.220 2.700 ;
        RECT 2579.940 1.820 2583.820 2.700 ;
        RECT 2585.540 1.820 2589.420 2.700 ;
        RECT 2591.140 1.820 2595.020 2.700 ;
        RECT 2596.740 1.820 2600.620 2.700 ;
        RECT 2602.340 1.820 2606.220 2.700 ;
        RECT 2607.940 1.820 2611.820 2.700 ;
        RECT 2613.540 1.820 2617.420 2.700 ;
        RECT 2619.140 1.820 2623.020 2.700 ;
        RECT 2624.740 1.820 2628.620 2.700 ;
        RECT 2630.340 1.820 2634.220 2.700 ;
        RECT 2635.940 1.820 2639.820 2.700 ;
        RECT 2641.540 1.820 2645.420 2.700 ;
        RECT 2647.140 1.820 2651.020 2.700 ;
        RECT 2652.740 1.820 2656.620 2.700 ;
        RECT 2658.340 1.820 2662.220 2.700 ;
        RECT 2663.940 1.820 2667.820 2.700 ;
        RECT 2669.540 1.820 2673.420 2.700 ;
        RECT 2675.140 1.820 2679.020 2.700 ;
        RECT 2680.740 1.820 2684.620 2.700 ;
        RECT 2686.340 1.820 2690.220 2.700 ;
        RECT 2691.940 1.820 2695.820 2.700 ;
        RECT 2697.540 1.820 2701.420 2.700 ;
        RECT 2703.140 1.820 2707.020 2.700 ;
        RECT 2708.740 1.820 2712.620 2.700 ;
        RECT 2714.340 1.820 2718.220 2.700 ;
        RECT 2719.940 1.820 2723.820 2.700 ;
        RECT 2725.540 1.820 2729.420 2.700 ;
        RECT 2731.140 1.820 2735.020 2.700 ;
        RECT 2736.740 1.820 2740.620 2.700 ;
        RECT 2742.340 1.820 2746.220 2.700 ;
        RECT 2747.940 1.820 2751.820 2.700 ;
        RECT 2753.540 1.820 2757.420 2.700 ;
        RECT 2759.140 1.820 2763.020 2.700 ;
        RECT 2764.740 1.820 2768.620 2.700 ;
        RECT 2770.340 1.820 2774.220 2.700 ;
        RECT 2775.940 1.820 2779.820 2.700 ;
        RECT 2781.540 1.820 2785.420 2.700 ;
        RECT 2787.140 1.820 2791.020 2.700 ;
        RECT 2792.740 1.820 2796.620 2.700 ;
        RECT 2798.340 1.820 2802.220 2.700 ;
        RECT 2803.940 1.820 2807.820 2.700 ;
        RECT 2809.540 1.820 2813.420 2.700 ;
        RECT 2815.140 1.820 2819.020 2.700 ;
        RECT 2820.740 1.820 2824.620 2.700 ;
        RECT 2826.340 1.820 2830.220 2.700 ;
        RECT 2831.940 1.820 2835.820 2.700 ;
        RECT 2837.540 1.820 2841.420 2.700 ;
        RECT 2843.140 1.820 2847.020 2.700 ;
        RECT 2848.740 1.820 2852.620 2.700 ;
        RECT 2854.340 1.820 2858.220 2.700 ;
        RECT 2859.940 1.820 2863.820 2.700 ;
        RECT 2865.540 1.820 2869.420 2.700 ;
        RECT 2871.140 1.820 2970.100 2.700 ;
      LAYER Metal3 ;
        RECT 1.820 2946.740 2978.500 2956.660 ;
        RECT 1.820 2945.060 2977.500 2946.740 ;
        RECT 2.700 2945.020 2977.500 2945.060 ;
        RECT 2.700 2943.340 2978.500 2945.020 ;
        RECT 1.820 2890.740 2978.500 2943.340 ;
        RECT 1.820 2890.180 2977.500 2890.740 ;
        RECT 2.700 2889.020 2977.500 2890.180 ;
        RECT 2.700 2888.460 2978.500 2889.020 ;
        RECT 1.820 2835.300 2978.500 2888.460 ;
        RECT 2.700 2834.740 2978.500 2835.300 ;
        RECT 2.700 2833.580 2977.500 2834.740 ;
        RECT 1.820 2833.020 2977.500 2833.580 ;
        RECT 1.820 2780.420 2978.500 2833.020 ;
        RECT 2.700 2778.740 2978.500 2780.420 ;
        RECT 2.700 2778.700 2977.500 2778.740 ;
        RECT 1.820 2777.020 2977.500 2778.700 ;
        RECT 1.820 2725.540 2978.500 2777.020 ;
        RECT 2.700 2723.820 2978.500 2725.540 ;
        RECT 1.820 2722.740 2978.500 2723.820 ;
        RECT 1.820 2721.020 2977.500 2722.740 ;
        RECT 1.820 2670.660 2978.500 2721.020 ;
        RECT 2.700 2668.940 2978.500 2670.660 ;
        RECT 1.820 2666.740 2978.500 2668.940 ;
        RECT 1.820 2665.020 2977.500 2666.740 ;
        RECT 1.820 2615.780 2978.500 2665.020 ;
        RECT 2.700 2614.060 2978.500 2615.780 ;
        RECT 1.820 2610.740 2978.500 2614.060 ;
        RECT 1.820 2609.020 2977.500 2610.740 ;
        RECT 1.820 2560.900 2978.500 2609.020 ;
        RECT 2.700 2559.180 2978.500 2560.900 ;
        RECT 1.820 2554.740 2978.500 2559.180 ;
        RECT 1.820 2553.020 2977.500 2554.740 ;
        RECT 1.820 2506.020 2978.500 2553.020 ;
        RECT 2.700 2504.300 2978.500 2506.020 ;
        RECT 1.820 2498.740 2978.500 2504.300 ;
        RECT 1.820 2497.020 2977.500 2498.740 ;
        RECT 1.820 2451.140 2978.500 2497.020 ;
        RECT 2.700 2449.420 2978.500 2451.140 ;
        RECT 1.820 2442.740 2978.500 2449.420 ;
        RECT 1.820 2441.020 2977.500 2442.740 ;
        RECT 1.820 2396.260 2978.500 2441.020 ;
        RECT 2.700 2394.540 2978.500 2396.260 ;
        RECT 1.820 2386.740 2978.500 2394.540 ;
        RECT 1.820 2385.020 2977.500 2386.740 ;
        RECT 1.820 2341.380 2978.500 2385.020 ;
        RECT 2.700 2339.660 2978.500 2341.380 ;
        RECT 1.820 2330.740 2978.500 2339.660 ;
        RECT 1.820 2329.020 2977.500 2330.740 ;
        RECT 1.820 2286.500 2978.500 2329.020 ;
        RECT 2.700 2284.780 2978.500 2286.500 ;
        RECT 1.820 2274.740 2978.500 2284.780 ;
        RECT 1.820 2273.020 2977.500 2274.740 ;
        RECT 1.820 2231.620 2978.500 2273.020 ;
        RECT 2.700 2229.900 2978.500 2231.620 ;
        RECT 1.820 2218.740 2978.500 2229.900 ;
        RECT 1.820 2217.020 2977.500 2218.740 ;
        RECT 1.820 2176.740 2978.500 2217.020 ;
        RECT 2.700 2175.020 2978.500 2176.740 ;
        RECT 1.820 2162.740 2978.500 2175.020 ;
        RECT 1.820 2161.020 2977.500 2162.740 ;
        RECT 1.820 2121.860 2978.500 2161.020 ;
        RECT 2.700 2120.140 2978.500 2121.860 ;
        RECT 1.820 2106.740 2978.500 2120.140 ;
        RECT 1.820 2105.020 2977.500 2106.740 ;
        RECT 1.820 2066.980 2978.500 2105.020 ;
        RECT 2.700 2065.260 2978.500 2066.980 ;
        RECT 1.820 2050.740 2978.500 2065.260 ;
        RECT 1.820 2049.020 2977.500 2050.740 ;
        RECT 1.820 2012.100 2978.500 2049.020 ;
        RECT 2.700 2010.380 2978.500 2012.100 ;
        RECT 1.820 1994.740 2978.500 2010.380 ;
        RECT 1.820 1993.020 2977.500 1994.740 ;
        RECT 1.820 1957.220 2978.500 1993.020 ;
        RECT 2.700 1955.500 2978.500 1957.220 ;
        RECT 1.820 1938.740 2978.500 1955.500 ;
        RECT 1.820 1937.020 2977.500 1938.740 ;
        RECT 1.820 1902.340 2978.500 1937.020 ;
        RECT 2.700 1900.620 2978.500 1902.340 ;
        RECT 1.820 1882.740 2978.500 1900.620 ;
        RECT 1.820 1881.020 2977.500 1882.740 ;
        RECT 1.820 1847.460 2978.500 1881.020 ;
        RECT 2.700 1845.740 2978.500 1847.460 ;
        RECT 1.820 1826.740 2978.500 1845.740 ;
        RECT 1.820 1825.020 2977.500 1826.740 ;
        RECT 1.820 1792.580 2978.500 1825.020 ;
        RECT 2.700 1790.860 2978.500 1792.580 ;
        RECT 1.820 1770.740 2978.500 1790.860 ;
        RECT 1.820 1769.020 2977.500 1770.740 ;
        RECT 1.820 1737.700 2978.500 1769.020 ;
        RECT 2.700 1735.980 2978.500 1737.700 ;
        RECT 1.820 1714.740 2978.500 1735.980 ;
        RECT 1.820 1713.020 2977.500 1714.740 ;
        RECT 1.820 1682.820 2978.500 1713.020 ;
        RECT 2.700 1681.100 2978.500 1682.820 ;
        RECT 1.820 1658.740 2978.500 1681.100 ;
        RECT 1.820 1657.020 2977.500 1658.740 ;
        RECT 1.820 1627.940 2978.500 1657.020 ;
        RECT 2.700 1626.220 2978.500 1627.940 ;
        RECT 1.820 1602.740 2978.500 1626.220 ;
        RECT 1.820 1601.020 2977.500 1602.740 ;
        RECT 1.820 1573.060 2978.500 1601.020 ;
        RECT 2.700 1571.340 2978.500 1573.060 ;
        RECT 1.820 1546.740 2978.500 1571.340 ;
        RECT 1.820 1545.020 2977.500 1546.740 ;
        RECT 1.820 1518.180 2978.500 1545.020 ;
        RECT 2.700 1516.460 2978.500 1518.180 ;
        RECT 1.820 1490.740 2978.500 1516.460 ;
        RECT 1.820 1489.020 2977.500 1490.740 ;
        RECT 1.820 1463.300 2978.500 1489.020 ;
        RECT 2.700 1461.580 2978.500 1463.300 ;
        RECT 1.820 1434.740 2978.500 1461.580 ;
        RECT 1.820 1433.020 2977.500 1434.740 ;
        RECT 1.820 1408.420 2978.500 1433.020 ;
        RECT 2.700 1406.700 2978.500 1408.420 ;
        RECT 1.820 1378.740 2978.500 1406.700 ;
        RECT 1.820 1377.020 2977.500 1378.740 ;
        RECT 1.820 1353.540 2978.500 1377.020 ;
        RECT 2.700 1351.820 2978.500 1353.540 ;
        RECT 1.820 1322.740 2978.500 1351.820 ;
        RECT 1.820 1321.020 2977.500 1322.740 ;
        RECT 1.820 1298.660 2978.500 1321.020 ;
        RECT 2.700 1296.940 2978.500 1298.660 ;
        RECT 1.820 1266.740 2978.500 1296.940 ;
        RECT 1.820 1265.020 2977.500 1266.740 ;
        RECT 1.820 1243.780 2978.500 1265.020 ;
        RECT 2.700 1242.060 2978.500 1243.780 ;
        RECT 1.820 1210.740 2978.500 1242.060 ;
        RECT 1.820 1209.020 2977.500 1210.740 ;
        RECT 1.820 1188.900 2978.500 1209.020 ;
        RECT 2.700 1187.180 2978.500 1188.900 ;
        RECT 1.820 1154.740 2978.500 1187.180 ;
        RECT 1.820 1153.020 2977.500 1154.740 ;
        RECT 1.820 1134.020 2978.500 1153.020 ;
        RECT 2.700 1132.300 2978.500 1134.020 ;
        RECT 1.820 1098.740 2978.500 1132.300 ;
        RECT 1.820 1097.020 2977.500 1098.740 ;
        RECT 1.820 1079.140 2978.500 1097.020 ;
        RECT 2.700 1077.420 2978.500 1079.140 ;
        RECT 1.820 1042.740 2978.500 1077.420 ;
        RECT 1.820 1041.020 2977.500 1042.740 ;
        RECT 1.820 1024.260 2978.500 1041.020 ;
        RECT 2.700 1022.540 2978.500 1024.260 ;
        RECT 1.820 986.740 2978.500 1022.540 ;
        RECT 1.820 985.020 2977.500 986.740 ;
        RECT 1.820 969.380 2978.500 985.020 ;
        RECT 2.700 967.660 2978.500 969.380 ;
        RECT 1.820 930.740 2978.500 967.660 ;
        RECT 1.820 929.020 2977.500 930.740 ;
        RECT 1.820 914.500 2978.500 929.020 ;
        RECT 2.700 912.780 2978.500 914.500 ;
        RECT 1.820 874.740 2978.500 912.780 ;
        RECT 1.820 873.020 2977.500 874.740 ;
        RECT 1.820 859.620 2978.500 873.020 ;
        RECT 2.700 857.900 2978.500 859.620 ;
        RECT 1.820 818.740 2978.500 857.900 ;
        RECT 1.820 817.020 2977.500 818.740 ;
        RECT 1.820 804.740 2978.500 817.020 ;
        RECT 2.700 803.020 2978.500 804.740 ;
        RECT 1.820 762.740 2978.500 803.020 ;
        RECT 1.820 761.020 2977.500 762.740 ;
        RECT 1.820 749.860 2978.500 761.020 ;
        RECT 2.700 748.140 2978.500 749.860 ;
        RECT 1.820 706.740 2978.500 748.140 ;
        RECT 1.820 705.020 2977.500 706.740 ;
        RECT 1.820 694.980 2978.500 705.020 ;
        RECT 2.700 693.260 2978.500 694.980 ;
        RECT 1.820 650.740 2978.500 693.260 ;
        RECT 1.820 649.020 2977.500 650.740 ;
        RECT 1.820 640.100 2978.500 649.020 ;
        RECT 2.700 638.380 2978.500 640.100 ;
        RECT 1.820 594.740 2978.500 638.380 ;
        RECT 1.820 593.020 2977.500 594.740 ;
        RECT 1.820 585.220 2978.500 593.020 ;
        RECT 2.700 583.500 2978.500 585.220 ;
        RECT 1.820 538.740 2978.500 583.500 ;
        RECT 1.820 537.020 2977.500 538.740 ;
        RECT 1.820 530.340 2978.500 537.020 ;
        RECT 2.700 528.620 2978.500 530.340 ;
        RECT 1.820 482.740 2978.500 528.620 ;
        RECT 1.820 481.020 2977.500 482.740 ;
        RECT 1.820 475.460 2978.500 481.020 ;
        RECT 2.700 473.740 2978.500 475.460 ;
        RECT 1.820 426.740 2978.500 473.740 ;
        RECT 1.820 425.020 2977.500 426.740 ;
        RECT 1.820 420.580 2978.500 425.020 ;
        RECT 2.700 418.860 2978.500 420.580 ;
        RECT 1.820 370.740 2978.500 418.860 ;
        RECT 1.820 369.020 2977.500 370.740 ;
        RECT 1.820 365.700 2978.500 369.020 ;
        RECT 2.700 363.980 2978.500 365.700 ;
        RECT 1.820 314.740 2978.500 363.980 ;
        RECT 1.820 313.020 2977.500 314.740 ;
        RECT 1.820 310.820 2978.500 313.020 ;
        RECT 2.700 309.100 2978.500 310.820 ;
        RECT 1.820 258.740 2978.500 309.100 ;
        RECT 1.820 257.020 2977.500 258.740 ;
        RECT 1.820 255.940 2978.500 257.020 ;
        RECT 2.700 254.220 2978.500 255.940 ;
        RECT 1.820 202.740 2978.500 254.220 ;
        RECT 1.820 201.060 2977.500 202.740 ;
        RECT 2.700 201.020 2977.500 201.060 ;
        RECT 2.700 199.340 2978.500 201.020 ;
        RECT 1.820 146.740 2978.500 199.340 ;
        RECT 1.820 146.180 2977.500 146.740 ;
        RECT 2.700 145.020 2977.500 146.180 ;
        RECT 2.700 144.460 2978.500 145.020 ;
        RECT 1.820 91.300 2978.500 144.460 ;
        RECT 2.700 90.740 2978.500 91.300 ;
        RECT 2.700 89.580 2977.500 90.740 ;
        RECT 1.820 89.020 2977.500 89.580 ;
        RECT 1.820 36.420 2978.500 89.020 ;
        RECT 2.700 34.740 2978.500 36.420 ;
        RECT 2.700 34.700 2977.500 34.740 ;
        RECT 1.820 33.020 2977.500 34.700 ;
        RECT 1.820 18.060 2978.500 33.020 ;
      LAYER Metal4 ;
        RECT 369.740 19.690 375.470 2298.150 ;
        RECT 379.170 19.690 394.070 2298.150 ;
        RECT 397.770 19.690 465.470 2298.150 ;
        RECT 469.170 19.690 484.070 2298.150 ;
        RECT 487.770 19.690 555.470 2298.150 ;
        RECT 559.170 19.690 574.070 2298.150 ;
        RECT 577.770 19.690 645.470 2298.150 ;
        RECT 649.170 19.690 664.070 2298.150 ;
        RECT 667.770 19.690 735.470 2298.150 ;
        RECT 739.170 19.690 754.070 2298.150 ;
        RECT 757.770 19.690 825.470 2298.150 ;
        RECT 829.170 19.690 844.070 2298.150 ;
        RECT 847.770 19.690 915.470 2298.150 ;
        RECT 919.170 19.690 934.070 2298.150 ;
        RECT 937.770 19.690 1005.470 2298.150 ;
        RECT 1009.170 19.690 1024.070 2298.150 ;
        RECT 1027.770 19.690 1095.470 2298.150 ;
        RECT 1099.170 19.690 1114.070 2298.150 ;
        RECT 1117.770 19.690 1185.470 2298.150 ;
        RECT 1189.170 19.690 1204.070 2298.150 ;
        RECT 1207.770 2284.360 1275.470 2298.150 ;
        RECT 1279.170 2284.360 1294.070 2298.150 ;
        RECT 1207.770 1695.400 1294.070 2284.360 ;
        RECT 1207.770 19.690 1275.470 1695.400 ;
        RECT 1279.170 19.690 1294.070 1695.400 ;
        RECT 1297.770 19.690 1365.470 2298.150 ;
        RECT 1369.170 19.690 1384.070 2298.150 ;
        RECT 1387.770 19.690 1455.470 2298.150 ;
        RECT 1459.170 19.690 1474.070 2298.150 ;
        RECT 1477.770 19.690 1545.470 2298.150 ;
        RECT 1549.170 19.690 1564.070 2298.150 ;
        RECT 1567.770 19.690 1635.470 2298.150 ;
        RECT 1639.170 19.690 1654.070 2298.150 ;
        RECT 1657.770 2280.610 1725.470 2298.150 ;
        RECT 1729.170 2280.610 1744.070 2298.150 ;
        RECT 1747.770 2280.610 1815.470 2298.150 ;
        RECT 1657.770 2247.950 1815.470 2280.610 ;
        RECT 1657.770 19.690 1725.470 2247.950 ;
        RECT 1729.170 19.690 1744.070 2247.950 ;
        RECT 1747.770 19.690 1815.470 2247.950 ;
        RECT 1819.170 19.690 1834.070 2298.150 ;
        RECT 1837.770 19.690 1905.470 2298.150 ;
        RECT 1909.170 19.690 1924.070 2298.150 ;
        RECT 1927.770 19.690 1995.470 2298.150 ;
        RECT 1999.170 19.690 2014.070 2298.150 ;
        RECT 2017.770 19.690 2085.470 2298.150 ;
        RECT 2089.170 19.690 2104.070 2298.150 ;
        RECT 2107.770 19.690 2175.470 2298.150 ;
        RECT 2179.170 19.690 2194.070 2298.150 ;
        RECT 2197.770 19.690 2265.470 2298.150 ;
        RECT 2269.170 19.690 2284.070 2298.150 ;
        RECT 2287.770 19.690 2355.470 2298.150 ;
        RECT 2359.170 19.690 2374.070 2298.150 ;
        RECT 2377.770 19.690 2445.470 2298.150 ;
        RECT 2449.170 19.690 2464.070 2298.150 ;
        RECT 2467.770 19.690 2513.140 2298.150 ;
  END
END user_project_wrapper
END LIBRARY

